module chacha20_serial_encoder (
    clear,
    reset,
    clock,
    set_state,
    round_input,
    round_output
);

    input clear;
    input reset;
    input clock;
    input set_state;
    input [511:0] round_input;
    output [511:0] round_output;

    /* signal declarations */
    wire vdd = 1'b1;
    wire [511:0] _17 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire _2;
    wire [511:0] _16 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire _4;
    wire _6;
    wire [383:0] _24;
    wire [31:0] _22 = 32'b00000000000000000000000000000001;
    wire [31:0] _21;
    wire [31:0] _23;
    wire [95:0] _20;
    wire [511:0] _25;
    wire _14 = 1'b1;
    wire _8;
    wire _15;
    wire [511:0] _26;
    wire [511:0] _9;
    reg [511:0] _19;
    wire [511:0] _28;
    wire [511:0] _10;
    wire [511:0] _12;
    wire [511:0] _29;

    /* logic */
    assign _2 = clear;
    assign _4 = reset;
    assign _6 = clock;
    assign _24 = _19[383:0];
    assign _21 = _19[415:384];
    assign _23 = _21 + _22;
    assign _20 = _19[511:416];
    assign _25 = { _20, _23, _24 };
    assign _8 = set_state;
    assign _15 = _8 == _14;
    assign _26 = _15 ? _12 : _25;
    assign _9 = _26;
    always @(posedge _6 or posedge _4) begin
        if (_4)
            _19 <= _16;
        else
            if (_2)
                _19 <= _17;
            else
                _19 <= _9;
    end
    chacha20_block
        _0
        ( .round_input(_19), .round_output(_28[511:0]) );
    assign _10 = _28;
    assign _12 = round_input;
    assign _29 = _12 ^ _10;

    /* aliases */

    /* output assignments */
    assign round_output = _29;

endmodule
