module poly1305_block (
    number_of_input_bytes_minus_one,
    round_input,
    accumulator,
    r,
    new_accumulator
);

    input [3:0] number_of_input_bytes_minus_one;
    input [127:0] round_input;
    input [129:0] accumulator;
    input [127:0] r;
    output [129:0] new_accumulator;

    /* signal declarations */
    wire [258:0] _49 = 259'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011;
    wire [258:0] _43;
    wire [257:0] _44;
    wire _42 = 1'b0;
    wire [258:0] _45;
    wire [258:0] _37 = 259'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101;
    wire [517:0] _38;
    wire [258:0] _39;
    wire [258:0] _36 = 259'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [517:0] _40;
    wire [258:0] _41;
    wire [258:0] _46;
    wire [129:0] _47;
    wire [128:0] _35 = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [258:0] _48;
    wire [517:0] _50;
    wire [258:0] _51;
    wire [129:0] _29 = 130'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _28 = 130'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _27 = 130'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _26 = 130'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _25 = 130'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _24 = 130'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _23 = 130'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _22 = 130'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _21 = 130'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _20 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
    wire [129:0] _19 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
    wire [129:0] _18 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
    wire [129:0] _17 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;
    wire [129:0] _16 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
    wire [129:0] _15 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
    wire [129:0] _14 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
    wire [3:0] _2;
    reg [129:0] _30;
    wire [127:0] _4;
    wire [1:0] _12 = 2'b00;
    wire [129:0] _13;
    wire [129:0] _31;
    wire [130:0] _32;
    wire [129:0] _6;
    wire gnd = 1'b0;
    wire [130:0] _11;
    wire [130:0] _33;
    wire [127:0] _8;
    wire [258:0] _34;
    wire [258:0] _52;
    wire [129:0] _53;

    /* logic */
    assign _43 = _34 - _41;
    assign _44 = _43[258:1];
    assign _45 = { _42, _44 };
    assign _38 = _34 * _37;
    assign _39 = _38[517:259];
    assign _40 = { _36, _39 };
    assign _41 = _40[258:0];
    assign _46 = _41 + _45;
    assign _47 = _46[258:129];
    assign _48 = { _35, _47 };
    assign _50 = _48 * _49;
    assign _51 = _50[258:0];
    assign _2 = number_of_input_bytes_minus_one;
    always @* begin
        case (_2)
        0: _30 <= _14;
        1: _30 <= _15;
        2: _30 <= _16;
        3: _30 <= _17;
        4: _30 <= _18;
        5: _30 <= _19;
        6: _30 <= _20;
        7: _30 <= _21;
        8: _30 <= _22;
        9: _30 <= _23;
        10: _30 <= _24;
        11: _30 <= _25;
        12: _30 <= _26;
        13: _30 <= _27;
        14: _30 <= _28;
        default: _30 <= _29;
        endcase
    end
    assign _4 = round_input;
    assign _13 = { _12, _4 };
    assign _31 = _13 | _30;
    assign _32 = { gnd, _31 };
    assign _6 = accumulator;
    assign _11 = { gnd, _6 };
    assign _33 = _11 + _32;
    assign _8 = r;
    assign _34 = _8 * _33;
    assign _52 = _34 - _51;
    assign _53 = _52[129:0];

    /* aliases */

    /* output assignments */
    assign new_accumulator = _53;

endmodule
