module chacha20_block_function_without_mixing (
    round_input,
    clear,
    clock,
    start,
    finished,
    round_output
);

    input [511:0] round_input;
    input clear;
    input clock;
    input start;
    output finished;
    output [511:0] round_output;

    /* signal declarations */
    wire [511:0] _26 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _25 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _2;
    wire [511:0] _23 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _24;
    wire [511:0] _28;
    wire [511:0] _3;
    wire [511:0] _30;
    wire [511:0] _4;
    wire [511:0] _31;
    wire [511:0] _32;
    wire [511:0] _5;
    reg [511:0] _27;
    wire [4:0] _38 = 5'b00000;
    wire vdd = 1'b1;
    wire [4:0] _17 = 5'b00000;
    wire _8;
    wire [4:0] _16 = 5'b00000;
    wire _10;
    wire [4:0] _35 = 5'b00001;
    wire [4:0] _36;
    wire [4:0] _33 = 5'b01001;
    wire _21 = 1'b1;
    wire _12;
    wire _22;
    wire [4:0] _34;
    wire [4:0] _15 = 5'b00000;
    wire _20;
    wire [4:0] _37;
    wire [4:0] _13;
    reg [4:0] _19;
    wire _39;

    /* logic */
    assign _2 = round_input;
    assign _24 = _22 ? _2 : _23;
    assign _28 = _20 ? _27 : _24;
    assign _3 = _28;
    chacha20_column_and_diagonal_round
        column_and_diagonal
        ( .round_input(_3), .round_output(_30[511:0]) );
    assign _4 = _30;
    assign _31 = _22 ? _4 : _27;
    assign _32 = _20 ? _4 : _31;
    assign _5 = _32;
    always @(posedge _10) begin
        if (_8)
            _27 <= _26;
        else
            _27 <= _5;
    end
    assign _8 = clear;
    assign _10 = clock;
    assign _36 = _19 - _35;
    assign _12 = start;
    assign _22 = _12 == _21;
    assign _34 = _22 ? _33 : _19;
    assign _20 = _15 < _19;
    assign _37 = _20 ? _36 : _34;
    assign _13 = _37;
    always @(posedge _10) begin
        if (_8)
            _19 <= _17;
        else
            _19 <= _13;
    end
    assign _39 = _19 == _38;

    /* aliases */

    /* output assignments */
    assign finished = _39;
    assign round_output = _27;

endmodule
