module chacha20_serial_encoder (
    clear,
    clock,
    set_state,
    round_input,
    round_output
);

    input clear;
    input clock;
    input set_state;
    input [511:0] round_input;
    output [511:0] round_output;

    /* signal declarations */
    wire [31:0] _2910;
    wire [31:0] _2909;
    wire [31:0] _2911;
    wire [31:0] _2907;
    wire [31:0] _2906;
    wire [31:0] _2908;
    wire [31:0] _2904;
    wire [31:0] _2903;
    wire [31:0] _2905;
    wire [31:0] _2901;
    wire [31:0] _2900;
    wire [31:0] _2902;
    wire [31:0] _2898;
    wire [31:0] _2897;
    wire [31:0] _2899;
    wire [31:0] _2895;
    wire [31:0] _2894;
    wire [31:0] _2896;
    wire [31:0] _2892;
    wire [31:0] _2891;
    wire [31:0] _2893;
    wire [31:0] _2889;
    wire [31:0] _2888;
    wire [31:0] _2890;
    wire [31:0] _2886;
    wire [31:0] _2885;
    wire [31:0] _2887;
    wire [31:0] _2883;
    wire [31:0] _2882;
    wire [31:0] _2884;
    wire [31:0] _2880;
    wire [31:0] _2879;
    wire [31:0] _2881;
    wire [31:0] _2877;
    wire [31:0] _2876;
    wire [31:0] _2878;
    wire [31:0] _2874;
    wire [31:0] _2873;
    wire [31:0] _2875;
    wire [31:0] _2871;
    wire [31:0] _2870;
    wire [31:0] _2872;
    wire [31:0] _2868;
    wire [31:0] _2867;
    wire [31:0] _2869;
    wire [447:0] _2863;
    wire [287:0] _2860;
    wire [127:0] _2857;
    wire [6:0] _2855;
    wire [7:0] _2850;
    wire [31:0] _2848;
    wire [23:0] _2849;
    wire [31:0] _2851;
    wire [31:0] _2852;
    wire [31:0] _2853;
    wire [24:0] _2854;
    wire [31:0] _2856;
    wire [95:0] _2845;
    wire [11:0] _2842;
    wire [15:0] _2837;
    wire [31:0] _2834;
    wire [31:0] _2835;
    wire [15:0] _2836;
    wire [31:0] _2838;
    wire [31:0] _2833;
    wire [31:0] _2839;
    wire [31:0] _2840;
    wire [19:0] _2841;
    wire [31:0] _2843;
    wire [31:0] _2831;
    wire [31:0] _2830;
    wire [31:0] _2832;
    wire [31:0] _2844;
    wire [415:0] _2827;
    wire [255:0] _2824;
    wire [223:0] _2821;
    wire [6:0] _2819;
    wire [7:0] _2814;
    wire [31:0] _2812;
    wire [23:0] _2813;
    wire [31:0] _2815;
    wire [31:0] _2816;
    wire [31:0] _2817;
    wire [24:0] _2818;
    wire [31:0] _2820;
    wire [63:0] _2809;
    wire [11:0] _2806;
    wire [15:0] _2801;
    wire [31:0] _2798;
    wire [31:0] _2799;
    wire [15:0] _2800;
    wire [31:0] _2802;
    wire [31:0] _2797;
    wire [31:0] _2803;
    wire [31:0] _2804;
    wire [19:0] _2805;
    wire [31:0] _2807;
    wire [31:0] _2795;
    wire [31:0] _2794;
    wire [31:0] _2796;
    wire [31:0] _2808;
    wire [383:0] _2791;
    wire [351:0] _2788;
    wire [191:0] _2785;
    wire [6:0] _2783;
    wire [7:0] _2778;
    wire [31:0] _2776;
    wire [23:0] _2777;
    wire [31:0] _2779;
    wire [31:0] _2780;
    wire [31:0] _2781;
    wire [24:0] _2782;
    wire [31:0] _2784;
    wire [31:0] _2773;
    wire [11:0] _2770;
    wire [15:0] _2765;
    wire [31:0] _2762;
    wire [31:0] _2763;
    wire [15:0] _2764;
    wire [31:0] _2766;
    wire [31:0] _2761;
    wire [31:0] _2767;
    wire [31:0] _2768;
    wire [19:0] _2769;
    wire [31:0] _2771;
    wire [31:0] _2759;
    wire [31:0] _2758;
    wire [31:0] _2760;
    wire [31:0] _2772;
    wire [319:0] _2753;
    wire [159:0] _2750;
    wire [6:0] _2748;
    wire [31:0] _2745;
    wire [31:0] _2746;
    wire [24:0] _2747;
    wire [31:0] _2749;
    wire [479:0] _2742;
    wire [511:0] _2743;
    wire [319:0] _2744;
    wire [511:0] _2751;
    wire [159:0] _2752;
    wire [511:0] _2754;
    wire [479:0] _2755;
    wire [7:0] _2740;
    wire [11:0] _2735;
    wire [31:0] _2731;
    wire [31:0] _2732;
    wire [31:0] _2733;
    wire [19:0] _2734;
    wire [31:0] _2736;
    wire [31:0] _2737;
    wire [15:0] _2729;
    wire [31:0] _2725;
    wire [31:0] _2724;
    wire [31:0] _2726;
    wire [351:0] _2719;
    wire [223:0] _2716;
    wire [6:0] _2714;
    wire [31:0] _2711;
    wire [31:0] _2712;
    wire [24:0] _2713;
    wire [31:0] _2715;
    wire [95:0] _2708;
    wire [383:0] _2707;
    wire [511:0] _2709;
    wire [255:0] _2710;
    wire [511:0] _2717;
    wire [127:0] _2718;
    wire [511:0] _2720;
    wire [479:0] _2721;
    wire [7:0] _2705;
    wire [11:0] _2700;
    wire [31:0] _2696;
    wire [31:0] _2697;
    wire [31:0] _2698;
    wire [19:0] _2699;
    wire [31:0] _2701;
    wire [31:0] _2702;
    wire [15:0] _2694;
    wire [31:0] _2690;
    wire [31:0] _2689;
    wire [31:0] _2691;
    wire [447:0] _2686;
    wire [319:0] _2683;
    wire [191:0] _2680;
    wire [6:0] _2678;
    wire [7:0] _2673;
    wire [31:0] _2671;
    wire [23:0] _2672;
    wire [31:0] _2674;
    wire [31:0] _2675;
    wire [31:0] _2676;
    wire [24:0] _2677;
    wire [31:0] _2679;
    wire [63:0] _2668;
    wire [11:0] _2665;
    wire [15:0] _2660;
    wire [31:0] _2657;
    wire [31:0] _2658;
    wire [15:0] _2659;
    wire [31:0] _2661;
    wire [31:0] _2656;
    wire [31:0] _2662;
    wire [31:0] _2663;
    wire [19:0] _2664;
    wire [31:0] _2666;
    wire [31:0] _2654;
    wire [31:0] _2653;
    wire [31:0] _2655;
    wire [31:0] _2667;
    wire [415:0] _2650;
    wire [287:0] _2647;
    wire [159:0] _2644;
    wire [6:0] _2642;
    wire [7:0] _2637;
    wire [31:0] _2635;
    wire [23:0] _2636;
    wire [31:0] _2638;
    wire [31:0] _2639;
    wire [31:0] _2640;
    wire [24:0] _2641;
    wire [31:0] _2643;
    wire [31:0] _2632;
    wire [11:0] _2629;
    wire [15:0] _2624;
    wire [31:0] _2621;
    wire [31:0] _2622;
    wire [15:0] _2623;
    wire [31:0] _2625;
    wire [31:0] _2620;
    wire [31:0] _2626;
    wire [31:0] _2627;
    wire [19:0] _2628;
    wire [31:0] _2630;
    wire [31:0] _2618;
    wire [31:0] _2617;
    wire [31:0] _2619;
    wire [31:0] _2631;
    wire [383:0] _2614;
    wire [255:0] _2611;
    wire [127:0] _2608;
    wire [6:0] _2606;
    wire [7:0] _2601;
    wire [31:0] _2599;
    wire [23:0] _2600;
    wire [31:0] _2602;
    wire [31:0] _2603;
    wire [31:0] _2604;
    wire [24:0] _2605;
    wire [31:0] _2607;
    wire [11:0] _2594;
    wire [15:0] _2589;
    wire [31:0] _2586;
    wire [31:0] _2587;
    wire [15:0] _2588;
    wire [31:0] _2590;
    wire [31:0] _2585;
    wire [31:0] _2591;
    wire [31:0] _2592;
    wire [19:0] _2593;
    wire [31:0] _2595;
    wire [31:0] _2583;
    wire [31:0] _2582;
    wire [31:0] _2584;
    wire [31:0] _2596;
    wire [447:0] _2579;
    wire [287:0] _2576;
    wire [127:0] _2573;
    wire [6:0] _2571;
    wire [7:0] _2566;
    wire [31:0] _2564;
    wire [23:0] _2565;
    wire [31:0] _2567;
    wire [31:0] _2568;
    wire [31:0] _2569;
    wire [24:0] _2570;
    wire [31:0] _2572;
    wire [95:0] _2561;
    wire [11:0] _2558;
    wire [15:0] _2553;
    wire [31:0] _2550;
    wire [31:0] _2551;
    wire [15:0] _2552;
    wire [31:0] _2554;
    wire [31:0] _2549;
    wire [31:0] _2555;
    wire [31:0] _2556;
    wire [19:0] _2557;
    wire [31:0] _2559;
    wire [31:0] _2547;
    wire [31:0] _2546;
    wire [31:0] _2548;
    wire [31:0] _2560;
    wire [415:0] _2543;
    wire [255:0] _2540;
    wire [223:0] _2537;
    wire [6:0] _2535;
    wire [7:0] _2530;
    wire [31:0] _2528;
    wire [23:0] _2529;
    wire [31:0] _2531;
    wire [31:0] _2532;
    wire [31:0] _2533;
    wire [24:0] _2534;
    wire [31:0] _2536;
    wire [63:0] _2525;
    wire [11:0] _2522;
    wire [15:0] _2517;
    wire [31:0] _2514;
    wire [31:0] _2515;
    wire [15:0] _2516;
    wire [31:0] _2518;
    wire [31:0] _2513;
    wire [31:0] _2519;
    wire [31:0] _2520;
    wire [19:0] _2521;
    wire [31:0] _2523;
    wire [31:0] _2511;
    wire [31:0] _2510;
    wire [31:0] _2512;
    wire [31:0] _2524;
    wire [383:0] _2507;
    wire [351:0] _2504;
    wire [191:0] _2501;
    wire [6:0] _2499;
    wire [7:0] _2494;
    wire [31:0] _2492;
    wire [23:0] _2493;
    wire [31:0] _2495;
    wire [31:0] _2496;
    wire [31:0] _2497;
    wire [24:0] _2498;
    wire [31:0] _2500;
    wire [31:0] _2489;
    wire [11:0] _2486;
    wire [15:0] _2481;
    wire [31:0] _2478;
    wire [31:0] _2479;
    wire [15:0] _2480;
    wire [31:0] _2482;
    wire [31:0] _2477;
    wire [31:0] _2483;
    wire [31:0] _2484;
    wire [19:0] _2485;
    wire [31:0] _2487;
    wire [31:0] _2475;
    wire [31:0] _2474;
    wire [31:0] _2476;
    wire [31:0] _2488;
    wire [319:0] _2469;
    wire [159:0] _2466;
    wire [6:0] _2464;
    wire [31:0] _2461;
    wire [31:0] _2462;
    wire [24:0] _2463;
    wire [31:0] _2465;
    wire [479:0] _2458;
    wire [511:0] _2459;
    wire [319:0] _2460;
    wire [511:0] _2467;
    wire [159:0] _2468;
    wire [511:0] _2470;
    wire [479:0] _2471;
    wire [7:0] _2456;
    wire [11:0] _2451;
    wire [31:0] _2447;
    wire [31:0] _2448;
    wire [31:0] _2449;
    wire [19:0] _2450;
    wire [31:0] _2452;
    wire [31:0] _2453;
    wire [15:0] _2445;
    wire [31:0] _2441;
    wire [31:0] _2440;
    wire [31:0] _2442;
    wire [351:0] _2435;
    wire [223:0] _2432;
    wire [6:0] _2430;
    wire [31:0] _2427;
    wire [31:0] _2428;
    wire [24:0] _2429;
    wire [31:0] _2431;
    wire [95:0] _2424;
    wire [383:0] _2423;
    wire [511:0] _2425;
    wire [255:0] _2426;
    wire [511:0] _2433;
    wire [127:0] _2434;
    wire [511:0] _2436;
    wire [479:0] _2437;
    wire [7:0] _2421;
    wire [11:0] _2416;
    wire [31:0] _2412;
    wire [31:0] _2413;
    wire [31:0] _2414;
    wire [19:0] _2415;
    wire [31:0] _2417;
    wire [31:0] _2418;
    wire [15:0] _2410;
    wire [31:0] _2406;
    wire [31:0] _2405;
    wire [31:0] _2407;
    wire [447:0] _2402;
    wire [319:0] _2399;
    wire [191:0] _2396;
    wire [6:0] _2394;
    wire [7:0] _2389;
    wire [31:0] _2387;
    wire [23:0] _2388;
    wire [31:0] _2390;
    wire [31:0] _2391;
    wire [31:0] _2392;
    wire [24:0] _2393;
    wire [31:0] _2395;
    wire [63:0] _2384;
    wire [11:0] _2381;
    wire [15:0] _2376;
    wire [31:0] _2373;
    wire [31:0] _2374;
    wire [15:0] _2375;
    wire [31:0] _2377;
    wire [31:0] _2372;
    wire [31:0] _2378;
    wire [31:0] _2379;
    wire [19:0] _2380;
    wire [31:0] _2382;
    wire [31:0] _2370;
    wire [31:0] _2369;
    wire [31:0] _2371;
    wire [31:0] _2383;
    wire [415:0] _2366;
    wire [287:0] _2363;
    wire [159:0] _2360;
    wire [6:0] _2358;
    wire [7:0] _2353;
    wire [31:0] _2351;
    wire [23:0] _2352;
    wire [31:0] _2354;
    wire [31:0] _2355;
    wire [31:0] _2356;
    wire [24:0] _2357;
    wire [31:0] _2359;
    wire [31:0] _2348;
    wire [11:0] _2345;
    wire [15:0] _2340;
    wire [31:0] _2337;
    wire [31:0] _2338;
    wire [15:0] _2339;
    wire [31:0] _2341;
    wire [31:0] _2336;
    wire [31:0] _2342;
    wire [31:0] _2343;
    wire [19:0] _2344;
    wire [31:0] _2346;
    wire [31:0] _2334;
    wire [31:0] _2333;
    wire [31:0] _2335;
    wire [31:0] _2347;
    wire [383:0] _2330;
    wire [255:0] _2327;
    wire [127:0] _2324;
    wire [6:0] _2322;
    wire [7:0] _2317;
    wire [31:0] _2315;
    wire [23:0] _2316;
    wire [31:0] _2318;
    wire [31:0] _2319;
    wire [31:0] _2320;
    wire [24:0] _2321;
    wire [31:0] _2323;
    wire [11:0] _2310;
    wire [15:0] _2305;
    wire [31:0] _2302;
    wire [31:0] _2303;
    wire [15:0] _2304;
    wire [31:0] _2306;
    wire [31:0] _2301;
    wire [31:0] _2307;
    wire [31:0] _2308;
    wire [19:0] _2309;
    wire [31:0] _2311;
    wire [31:0] _2299;
    wire [31:0] _2298;
    wire [31:0] _2300;
    wire [31:0] _2312;
    wire [447:0] _2295;
    wire [287:0] _2292;
    wire [127:0] _2289;
    wire [6:0] _2287;
    wire [7:0] _2282;
    wire [31:0] _2280;
    wire [23:0] _2281;
    wire [31:0] _2283;
    wire [31:0] _2284;
    wire [31:0] _2285;
    wire [24:0] _2286;
    wire [31:0] _2288;
    wire [95:0] _2277;
    wire [11:0] _2274;
    wire [15:0] _2269;
    wire [31:0] _2266;
    wire [31:0] _2267;
    wire [15:0] _2268;
    wire [31:0] _2270;
    wire [31:0] _2265;
    wire [31:0] _2271;
    wire [31:0] _2272;
    wire [19:0] _2273;
    wire [31:0] _2275;
    wire [31:0] _2263;
    wire [31:0] _2262;
    wire [31:0] _2264;
    wire [31:0] _2276;
    wire [415:0] _2259;
    wire [255:0] _2256;
    wire [223:0] _2253;
    wire [6:0] _2251;
    wire [7:0] _2246;
    wire [31:0] _2244;
    wire [23:0] _2245;
    wire [31:0] _2247;
    wire [31:0] _2248;
    wire [31:0] _2249;
    wire [24:0] _2250;
    wire [31:0] _2252;
    wire [63:0] _2241;
    wire [11:0] _2238;
    wire [15:0] _2233;
    wire [31:0] _2230;
    wire [31:0] _2231;
    wire [15:0] _2232;
    wire [31:0] _2234;
    wire [31:0] _2229;
    wire [31:0] _2235;
    wire [31:0] _2236;
    wire [19:0] _2237;
    wire [31:0] _2239;
    wire [31:0] _2227;
    wire [31:0] _2226;
    wire [31:0] _2228;
    wire [31:0] _2240;
    wire [383:0] _2223;
    wire [351:0] _2220;
    wire [191:0] _2217;
    wire [6:0] _2215;
    wire [7:0] _2210;
    wire [31:0] _2208;
    wire [23:0] _2209;
    wire [31:0] _2211;
    wire [31:0] _2212;
    wire [31:0] _2213;
    wire [24:0] _2214;
    wire [31:0] _2216;
    wire [31:0] _2205;
    wire [11:0] _2202;
    wire [15:0] _2197;
    wire [31:0] _2194;
    wire [31:0] _2195;
    wire [15:0] _2196;
    wire [31:0] _2198;
    wire [31:0] _2193;
    wire [31:0] _2199;
    wire [31:0] _2200;
    wire [19:0] _2201;
    wire [31:0] _2203;
    wire [31:0] _2191;
    wire [31:0] _2190;
    wire [31:0] _2192;
    wire [31:0] _2204;
    wire [319:0] _2185;
    wire [159:0] _2182;
    wire [6:0] _2180;
    wire [31:0] _2177;
    wire [31:0] _2178;
    wire [24:0] _2179;
    wire [31:0] _2181;
    wire [479:0] _2174;
    wire [511:0] _2175;
    wire [319:0] _2176;
    wire [511:0] _2183;
    wire [159:0] _2184;
    wire [511:0] _2186;
    wire [479:0] _2187;
    wire [7:0] _2172;
    wire [11:0] _2167;
    wire [31:0] _2163;
    wire [31:0] _2164;
    wire [31:0] _2165;
    wire [19:0] _2166;
    wire [31:0] _2168;
    wire [31:0] _2169;
    wire [15:0] _2161;
    wire [31:0] _2157;
    wire [31:0] _2156;
    wire [31:0] _2158;
    wire [351:0] _2151;
    wire [223:0] _2148;
    wire [6:0] _2146;
    wire [31:0] _2143;
    wire [31:0] _2144;
    wire [24:0] _2145;
    wire [31:0] _2147;
    wire [95:0] _2140;
    wire [383:0] _2139;
    wire [511:0] _2141;
    wire [255:0] _2142;
    wire [511:0] _2149;
    wire [127:0] _2150;
    wire [511:0] _2152;
    wire [479:0] _2153;
    wire [7:0] _2137;
    wire [11:0] _2132;
    wire [31:0] _2128;
    wire [31:0] _2129;
    wire [31:0] _2130;
    wire [19:0] _2131;
    wire [31:0] _2133;
    wire [31:0] _2134;
    wire [15:0] _2126;
    wire [31:0] _2122;
    wire [31:0] _2121;
    wire [31:0] _2123;
    wire [447:0] _2118;
    wire [319:0] _2115;
    wire [191:0] _2112;
    wire [6:0] _2110;
    wire [7:0] _2105;
    wire [31:0] _2103;
    wire [23:0] _2104;
    wire [31:0] _2106;
    wire [31:0] _2107;
    wire [31:0] _2108;
    wire [24:0] _2109;
    wire [31:0] _2111;
    wire [63:0] _2100;
    wire [11:0] _2097;
    wire [15:0] _2092;
    wire [31:0] _2089;
    wire [31:0] _2090;
    wire [15:0] _2091;
    wire [31:0] _2093;
    wire [31:0] _2088;
    wire [31:0] _2094;
    wire [31:0] _2095;
    wire [19:0] _2096;
    wire [31:0] _2098;
    wire [31:0] _2086;
    wire [31:0] _2085;
    wire [31:0] _2087;
    wire [31:0] _2099;
    wire [415:0] _2082;
    wire [287:0] _2079;
    wire [159:0] _2076;
    wire [6:0] _2074;
    wire [7:0] _2069;
    wire [31:0] _2067;
    wire [23:0] _2068;
    wire [31:0] _2070;
    wire [31:0] _2071;
    wire [31:0] _2072;
    wire [24:0] _2073;
    wire [31:0] _2075;
    wire [31:0] _2064;
    wire [11:0] _2061;
    wire [15:0] _2056;
    wire [31:0] _2053;
    wire [31:0] _2054;
    wire [15:0] _2055;
    wire [31:0] _2057;
    wire [31:0] _2052;
    wire [31:0] _2058;
    wire [31:0] _2059;
    wire [19:0] _2060;
    wire [31:0] _2062;
    wire [31:0] _2050;
    wire [31:0] _2049;
    wire [31:0] _2051;
    wire [31:0] _2063;
    wire [383:0] _2046;
    wire [255:0] _2043;
    wire [127:0] _2040;
    wire [6:0] _2038;
    wire [7:0] _2033;
    wire [31:0] _2031;
    wire [23:0] _2032;
    wire [31:0] _2034;
    wire [31:0] _2035;
    wire [31:0] _2036;
    wire [24:0] _2037;
    wire [31:0] _2039;
    wire [11:0] _2026;
    wire [15:0] _2021;
    wire [31:0] _2018;
    wire [31:0] _2019;
    wire [15:0] _2020;
    wire [31:0] _2022;
    wire [31:0] _2017;
    wire [31:0] _2023;
    wire [31:0] _2024;
    wire [19:0] _2025;
    wire [31:0] _2027;
    wire [31:0] _2015;
    wire [31:0] _2014;
    wire [31:0] _2016;
    wire [31:0] _2028;
    wire [447:0] _2011;
    wire [287:0] _2008;
    wire [127:0] _2005;
    wire [6:0] _2003;
    wire [7:0] _1998;
    wire [31:0] _1996;
    wire [23:0] _1997;
    wire [31:0] _1999;
    wire [31:0] _2000;
    wire [31:0] _2001;
    wire [24:0] _2002;
    wire [31:0] _2004;
    wire [95:0] _1993;
    wire [11:0] _1990;
    wire [15:0] _1985;
    wire [31:0] _1982;
    wire [31:0] _1983;
    wire [15:0] _1984;
    wire [31:0] _1986;
    wire [31:0] _1981;
    wire [31:0] _1987;
    wire [31:0] _1988;
    wire [19:0] _1989;
    wire [31:0] _1991;
    wire [31:0] _1979;
    wire [31:0] _1978;
    wire [31:0] _1980;
    wire [31:0] _1992;
    wire [415:0] _1975;
    wire [255:0] _1972;
    wire [223:0] _1969;
    wire [6:0] _1967;
    wire [7:0] _1962;
    wire [31:0] _1960;
    wire [23:0] _1961;
    wire [31:0] _1963;
    wire [31:0] _1964;
    wire [31:0] _1965;
    wire [24:0] _1966;
    wire [31:0] _1968;
    wire [63:0] _1957;
    wire [11:0] _1954;
    wire [15:0] _1949;
    wire [31:0] _1946;
    wire [31:0] _1947;
    wire [15:0] _1948;
    wire [31:0] _1950;
    wire [31:0] _1945;
    wire [31:0] _1951;
    wire [31:0] _1952;
    wire [19:0] _1953;
    wire [31:0] _1955;
    wire [31:0] _1943;
    wire [31:0] _1942;
    wire [31:0] _1944;
    wire [31:0] _1956;
    wire [383:0] _1939;
    wire [351:0] _1936;
    wire [191:0] _1933;
    wire [6:0] _1931;
    wire [7:0] _1926;
    wire [31:0] _1924;
    wire [23:0] _1925;
    wire [31:0] _1927;
    wire [31:0] _1928;
    wire [31:0] _1929;
    wire [24:0] _1930;
    wire [31:0] _1932;
    wire [31:0] _1921;
    wire [11:0] _1918;
    wire [15:0] _1913;
    wire [31:0] _1910;
    wire [31:0] _1911;
    wire [15:0] _1912;
    wire [31:0] _1914;
    wire [31:0] _1909;
    wire [31:0] _1915;
    wire [31:0] _1916;
    wire [19:0] _1917;
    wire [31:0] _1919;
    wire [31:0] _1907;
    wire [31:0] _1906;
    wire [31:0] _1908;
    wire [31:0] _1920;
    wire [319:0] _1901;
    wire [159:0] _1898;
    wire [6:0] _1896;
    wire [31:0] _1893;
    wire [31:0] _1894;
    wire [24:0] _1895;
    wire [31:0] _1897;
    wire [479:0] _1890;
    wire [511:0] _1891;
    wire [319:0] _1892;
    wire [511:0] _1899;
    wire [159:0] _1900;
    wire [511:0] _1902;
    wire [479:0] _1903;
    wire [7:0] _1888;
    wire [11:0] _1883;
    wire [31:0] _1879;
    wire [31:0] _1880;
    wire [31:0] _1881;
    wire [19:0] _1882;
    wire [31:0] _1884;
    wire [31:0] _1885;
    wire [15:0] _1877;
    wire [31:0] _1873;
    wire [31:0] _1872;
    wire [31:0] _1874;
    wire [351:0] _1867;
    wire [223:0] _1864;
    wire [6:0] _1862;
    wire [31:0] _1859;
    wire [31:0] _1860;
    wire [24:0] _1861;
    wire [31:0] _1863;
    wire [95:0] _1856;
    wire [383:0] _1855;
    wire [511:0] _1857;
    wire [255:0] _1858;
    wire [511:0] _1865;
    wire [127:0] _1866;
    wire [511:0] _1868;
    wire [479:0] _1869;
    wire [7:0] _1853;
    wire [11:0] _1848;
    wire [31:0] _1844;
    wire [31:0] _1845;
    wire [31:0] _1846;
    wire [19:0] _1847;
    wire [31:0] _1849;
    wire [31:0] _1850;
    wire [15:0] _1842;
    wire [31:0] _1838;
    wire [31:0] _1837;
    wire [31:0] _1839;
    wire [447:0] _1834;
    wire [319:0] _1831;
    wire [191:0] _1828;
    wire [6:0] _1826;
    wire [7:0] _1821;
    wire [31:0] _1819;
    wire [23:0] _1820;
    wire [31:0] _1822;
    wire [31:0] _1823;
    wire [31:0] _1824;
    wire [24:0] _1825;
    wire [31:0] _1827;
    wire [63:0] _1816;
    wire [11:0] _1813;
    wire [15:0] _1808;
    wire [31:0] _1805;
    wire [31:0] _1806;
    wire [15:0] _1807;
    wire [31:0] _1809;
    wire [31:0] _1804;
    wire [31:0] _1810;
    wire [31:0] _1811;
    wire [19:0] _1812;
    wire [31:0] _1814;
    wire [31:0] _1802;
    wire [31:0] _1801;
    wire [31:0] _1803;
    wire [31:0] _1815;
    wire [415:0] _1798;
    wire [287:0] _1795;
    wire [159:0] _1792;
    wire [6:0] _1790;
    wire [7:0] _1785;
    wire [31:0] _1783;
    wire [23:0] _1784;
    wire [31:0] _1786;
    wire [31:0] _1787;
    wire [31:0] _1788;
    wire [24:0] _1789;
    wire [31:0] _1791;
    wire [31:0] _1780;
    wire [11:0] _1777;
    wire [15:0] _1772;
    wire [31:0] _1769;
    wire [31:0] _1770;
    wire [15:0] _1771;
    wire [31:0] _1773;
    wire [31:0] _1768;
    wire [31:0] _1774;
    wire [31:0] _1775;
    wire [19:0] _1776;
    wire [31:0] _1778;
    wire [31:0] _1766;
    wire [31:0] _1765;
    wire [31:0] _1767;
    wire [31:0] _1779;
    wire [383:0] _1762;
    wire [255:0] _1759;
    wire [127:0] _1756;
    wire [6:0] _1754;
    wire [7:0] _1749;
    wire [31:0] _1747;
    wire [23:0] _1748;
    wire [31:0] _1750;
    wire [31:0] _1751;
    wire [31:0] _1752;
    wire [24:0] _1753;
    wire [31:0] _1755;
    wire [11:0] _1742;
    wire [15:0] _1737;
    wire [31:0] _1734;
    wire [31:0] _1735;
    wire [15:0] _1736;
    wire [31:0] _1738;
    wire [31:0] _1733;
    wire [31:0] _1739;
    wire [31:0] _1740;
    wire [19:0] _1741;
    wire [31:0] _1743;
    wire [31:0] _1731;
    wire [31:0] _1730;
    wire [31:0] _1732;
    wire [31:0] _1744;
    wire [447:0] _1727;
    wire [287:0] _1724;
    wire [127:0] _1721;
    wire [6:0] _1719;
    wire [7:0] _1714;
    wire [31:0] _1712;
    wire [23:0] _1713;
    wire [31:0] _1715;
    wire [31:0] _1716;
    wire [31:0] _1717;
    wire [24:0] _1718;
    wire [31:0] _1720;
    wire [95:0] _1709;
    wire [11:0] _1706;
    wire [15:0] _1701;
    wire [31:0] _1698;
    wire [31:0] _1699;
    wire [15:0] _1700;
    wire [31:0] _1702;
    wire [31:0] _1697;
    wire [31:0] _1703;
    wire [31:0] _1704;
    wire [19:0] _1705;
    wire [31:0] _1707;
    wire [31:0] _1695;
    wire [31:0] _1694;
    wire [31:0] _1696;
    wire [31:0] _1708;
    wire [415:0] _1691;
    wire [255:0] _1688;
    wire [223:0] _1685;
    wire [6:0] _1683;
    wire [7:0] _1678;
    wire [31:0] _1676;
    wire [23:0] _1677;
    wire [31:0] _1679;
    wire [31:0] _1680;
    wire [31:0] _1681;
    wire [24:0] _1682;
    wire [31:0] _1684;
    wire [63:0] _1673;
    wire [11:0] _1670;
    wire [15:0] _1665;
    wire [31:0] _1662;
    wire [31:0] _1663;
    wire [15:0] _1664;
    wire [31:0] _1666;
    wire [31:0] _1661;
    wire [31:0] _1667;
    wire [31:0] _1668;
    wire [19:0] _1669;
    wire [31:0] _1671;
    wire [31:0] _1659;
    wire [31:0] _1658;
    wire [31:0] _1660;
    wire [31:0] _1672;
    wire [383:0] _1655;
    wire [351:0] _1652;
    wire [191:0] _1649;
    wire [6:0] _1647;
    wire [7:0] _1642;
    wire [31:0] _1640;
    wire [23:0] _1641;
    wire [31:0] _1643;
    wire [31:0] _1644;
    wire [31:0] _1645;
    wire [24:0] _1646;
    wire [31:0] _1648;
    wire [31:0] _1637;
    wire [11:0] _1634;
    wire [15:0] _1629;
    wire [31:0] _1626;
    wire [31:0] _1627;
    wire [15:0] _1628;
    wire [31:0] _1630;
    wire [31:0] _1625;
    wire [31:0] _1631;
    wire [31:0] _1632;
    wire [19:0] _1633;
    wire [31:0] _1635;
    wire [31:0] _1623;
    wire [31:0] _1622;
    wire [31:0] _1624;
    wire [31:0] _1636;
    wire [319:0] _1617;
    wire [159:0] _1614;
    wire [6:0] _1612;
    wire [31:0] _1609;
    wire [31:0] _1610;
    wire [24:0] _1611;
    wire [31:0] _1613;
    wire [479:0] _1606;
    wire [511:0] _1607;
    wire [319:0] _1608;
    wire [511:0] _1615;
    wire [159:0] _1616;
    wire [511:0] _1618;
    wire [479:0] _1619;
    wire [7:0] _1604;
    wire [11:0] _1599;
    wire [31:0] _1595;
    wire [31:0] _1596;
    wire [31:0] _1597;
    wire [19:0] _1598;
    wire [31:0] _1600;
    wire [31:0] _1601;
    wire [15:0] _1593;
    wire [31:0] _1589;
    wire [31:0] _1588;
    wire [31:0] _1590;
    wire [351:0] _1583;
    wire [223:0] _1580;
    wire [6:0] _1578;
    wire [31:0] _1575;
    wire [31:0] _1576;
    wire [24:0] _1577;
    wire [31:0] _1579;
    wire [95:0] _1572;
    wire [383:0] _1571;
    wire [511:0] _1573;
    wire [255:0] _1574;
    wire [511:0] _1581;
    wire [127:0] _1582;
    wire [511:0] _1584;
    wire [479:0] _1585;
    wire [7:0] _1569;
    wire [11:0] _1564;
    wire [31:0] _1560;
    wire [31:0] _1561;
    wire [31:0] _1562;
    wire [19:0] _1563;
    wire [31:0] _1565;
    wire [31:0] _1566;
    wire [15:0] _1558;
    wire [31:0] _1554;
    wire [31:0] _1553;
    wire [31:0] _1555;
    wire [447:0] _1550;
    wire [319:0] _1547;
    wire [191:0] _1544;
    wire [6:0] _1542;
    wire [7:0] _1537;
    wire [31:0] _1535;
    wire [23:0] _1536;
    wire [31:0] _1538;
    wire [31:0] _1539;
    wire [31:0] _1540;
    wire [24:0] _1541;
    wire [31:0] _1543;
    wire [63:0] _1532;
    wire [11:0] _1529;
    wire [15:0] _1524;
    wire [31:0] _1521;
    wire [31:0] _1522;
    wire [15:0] _1523;
    wire [31:0] _1525;
    wire [31:0] _1520;
    wire [31:0] _1526;
    wire [31:0] _1527;
    wire [19:0] _1528;
    wire [31:0] _1530;
    wire [31:0] _1518;
    wire [31:0] _1517;
    wire [31:0] _1519;
    wire [31:0] _1531;
    wire [415:0] _1514;
    wire [287:0] _1511;
    wire [159:0] _1508;
    wire [6:0] _1506;
    wire [7:0] _1501;
    wire [31:0] _1499;
    wire [23:0] _1500;
    wire [31:0] _1502;
    wire [31:0] _1503;
    wire [31:0] _1504;
    wire [24:0] _1505;
    wire [31:0] _1507;
    wire [31:0] _1496;
    wire [11:0] _1493;
    wire [15:0] _1488;
    wire [31:0] _1485;
    wire [31:0] _1486;
    wire [15:0] _1487;
    wire [31:0] _1489;
    wire [31:0] _1484;
    wire [31:0] _1490;
    wire [31:0] _1491;
    wire [19:0] _1492;
    wire [31:0] _1494;
    wire [31:0] _1482;
    wire [31:0] _1481;
    wire [31:0] _1483;
    wire [31:0] _1495;
    wire [383:0] _1478;
    wire [255:0] _1475;
    wire [127:0] _1472;
    wire [6:0] _1470;
    wire [7:0] _1465;
    wire [31:0] _1463;
    wire [23:0] _1464;
    wire [31:0] _1466;
    wire [31:0] _1467;
    wire [31:0] _1468;
    wire [24:0] _1469;
    wire [31:0] _1471;
    wire [11:0] _1458;
    wire [15:0] _1453;
    wire [31:0] _1450;
    wire [31:0] _1451;
    wire [15:0] _1452;
    wire [31:0] _1454;
    wire [31:0] _1449;
    wire [31:0] _1455;
    wire [31:0] _1456;
    wire [19:0] _1457;
    wire [31:0] _1459;
    wire [31:0] _1447;
    wire [31:0] _1446;
    wire [31:0] _1448;
    wire [31:0] _1460;
    wire [447:0] _1443;
    wire [287:0] _1440;
    wire [127:0] _1437;
    wire [6:0] _1435;
    wire [7:0] _1430;
    wire [31:0] _1428;
    wire [23:0] _1429;
    wire [31:0] _1431;
    wire [31:0] _1432;
    wire [31:0] _1433;
    wire [24:0] _1434;
    wire [31:0] _1436;
    wire [95:0] _1425;
    wire [11:0] _1422;
    wire [15:0] _1417;
    wire [31:0] _1414;
    wire [31:0] _1415;
    wire [15:0] _1416;
    wire [31:0] _1418;
    wire [31:0] _1413;
    wire [31:0] _1419;
    wire [31:0] _1420;
    wire [19:0] _1421;
    wire [31:0] _1423;
    wire [31:0] _1411;
    wire [31:0] _1410;
    wire [31:0] _1412;
    wire [31:0] _1424;
    wire [415:0] _1407;
    wire [255:0] _1404;
    wire [223:0] _1401;
    wire [6:0] _1399;
    wire [7:0] _1394;
    wire [31:0] _1392;
    wire [23:0] _1393;
    wire [31:0] _1395;
    wire [31:0] _1396;
    wire [31:0] _1397;
    wire [24:0] _1398;
    wire [31:0] _1400;
    wire [63:0] _1389;
    wire [11:0] _1386;
    wire [15:0] _1381;
    wire [31:0] _1378;
    wire [31:0] _1379;
    wire [15:0] _1380;
    wire [31:0] _1382;
    wire [31:0] _1377;
    wire [31:0] _1383;
    wire [31:0] _1384;
    wire [19:0] _1385;
    wire [31:0] _1387;
    wire [31:0] _1375;
    wire [31:0] _1374;
    wire [31:0] _1376;
    wire [31:0] _1388;
    wire [383:0] _1371;
    wire [351:0] _1368;
    wire [191:0] _1365;
    wire [6:0] _1363;
    wire [7:0] _1358;
    wire [31:0] _1356;
    wire [23:0] _1357;
    wire [31:0] _1359;
    wire [31:0] _1360;
    wire [31:0] _1361;
    wire [24:0] _1362;
    wire [31:0] _1364;
    wire [31:0] _1353;
    wire [11:0] _1350;
    wire [15:0] _1345;
    wire [31:0] _1342;
    wire [31:0] _1343;
    wire [15:0] _1344;
    wire [31:0] _1346;
    wire [31:0] _1341;
    wire [31:0] _1347;
    wire [31:0] _1348;
    wire [19:0] _1349;
    wire [31:0] _1351;
    wire [31:0] _1339;
    wire [31:0] _1338;
    wire [31:0] _1340;
    wire [31:0] _1352;
    wire [319:0] _1333;
    wire [159:0] _1330;
    wire [6:0] _1328;
    wire [31:0] _1325;
    wire [31:0] _1326;
    wire [24:0] _1327;
    wire [31:0] _1329;
    wire [479:0] _1322;
    wire [511:0] _1323;
    wire [319:0] _1324;
    wire [511:0] _1331;
    wire [159:0] _1332;
    wire [511:0] _1334;
    wire [479:0] _1335;
    wire [7:0] _1320;
    wire [11:0] _1315;
    wire [31:0] _1311;
    wire [31:0] _1312;
    wire [31:0] _1313;
    wire [19:0] _1314;
    wire [31:0] _1316;
    wire [31:0] _1317;
    wire [15:0] _1309;
    wire [31:0] _1305;
    wire [31:0] _1304;
    wire [31:0] _1306;
    wire [351:0] _1299;
    wire [223:0] _1296;
    wire [6:0] _1294;
    wire [31:0] _1291;
    wire [31:0] _1292;
    wire [24:0] _1293;
    wire [31:0] _1295;
    wire [95:0] _1288;
    wire [383:0] _1287;
    wire [511:0] _1289;
    wire [255:0] _1290;
    wire [511:0] _1297;
    wire [127:0] _1298;
    wire [511:0] _1300;
    wire [479:0] _1301;
    wire [7:0] _1285;
    wire [11:0] _1280;
    wire [31:0] _1276;
    wire [31:0] _1277;
    wire [31:0] _1278;
    wire [19:0] _1279;
    wire [31:0] _1281;
    wire [31:0] _1282;
    wire [15:0] _1274;
    wire [31:0] _1270;
    wire [31:0] _1269;
    wire [31:0] _1271;
    wire [447:0] _1266;
    wire [319:0] _1263;
    wire [191:0] _1260;
    wire [6:0] _1258;
    wire [7:0] _1253;
    wire [31:0] _1251;
    wire [23:0] _1252;
    wire [31:0] _1254;
    wire [31:0] _1255;
    wire [31:0] _1256;
    wire [24:0] _1257;
    wire [31:0] _1259;
    wire [63:0] _1248;
    wire [11:0] _1245;
    wire [15:0] _1240;
    wire [31:0] _1237;
    wire [31:0] _1238;
    wire [15:0] _1239;
    wire [31:0] _1241;
    wire [31:0] _1236;
    wire [31:0] _1242;
    wire [31:0] _1243;
    wire [19:0] _1244;
    wire [31:0] _1246;
    wire [31:0] _1234;
    wire [31:0] _1233;
    wire [31:0] _1235;
    wire [31:0] _1247;
    wire [415:0] _1230;
    wire [287:0] _1227;
    wire [159:0] _1224;
    wire [6:0] _1222;
    wire [7:0] _1217;
    wire [31:0] _1215;
    wire [23:0] _1216;
    wire [31:0] _1218;
    wire [31:0] _1219;
    wire [31:0] _1220;
    wire [24:0] _1221;
    wire [31:0] _1223;
    wire [31:0] _1212;
    wire [11:0] _1209;
    wire [15:0] _1204;
    wire [31:0] _1201;
    wire [31:0] _1202;
    wire [15:0] _1203;
    wire [31:0] _1205;
    wire [31:0] _1200;
    wire [31:0] _1206;
    wire [31:0] _1207;
    wire [19:0] _1208;
    wire [31:0] _1210;
    wire [31:0] _1198;
    wire [31:0] _1197;
    wire [31:0] _1199;
    wire [31:0] _1211;
    wire [383:0] _1194;
    wire [255:0] _1191;
    wire [127:0] _1188;
    wire [6:0] _1186;
    wire [7:0] _1181;
    wire [31:0] _1179;
    wire [23:0] _1180;
    wire [31:0] _1182;
    wire [31:0] _1183;
    wire [31:0] _1184;
    wire [24:0] _1185;
    wire [31:0] _1187;
    wire [11:0] _1174;
    wire [15:0] _1169;
    wire [31:0] _1166;
    wire [31:0] _1167;
    wire [15:0] _1168;
    wire [31:0] _1170;
    wire [31:0] _1165;
    wire [31:0] _1171;
    wire [31:0] _1172;
    wire [19:0] _1173;
    wire [31:0] _1175;
    wire [31:0] _1163;
    wire [31:0] _1162;
    wire [31:0] _1164;
    wire [31:0] _1176;
    wire [447:0] _1159;
    wire [287:0] _1156;
    wire [127:0] _1153;
    wire [6:0] _1151;
    wire [7:0] _1146;
    wire [31:0] _1144;
    wire [23:0] _1145;
    wire [31:0] _1147;
    wire [31:0] _1148;
    wire [31:0] _1149;
    wire [24:0] _1150;
    wire [31:0] _1152;
    wire [95:0] _1141;
    wire [11:0] _1138;
    wire [15:0] _1133;
    wire [31:0] _1130;
    wire [31:0] _1131;
    wire [15:0] _1132;
    wire [31:0] _1134;
    wire [31:0] _1129;
    wire [31:0] _1135;
    wire [31:0] _1136;
    wire [19:0] _1137;
    wire [31:0] _1139;
    wire [31:0] _1127;
    wire [31:0] _1126;
    wire [31:0] _1128;
    wire [31:0] _1140;
    wire [415:0] _1123;
    wire [255:0] _1120;
    wire [223:0] _1117;
    wire [6:0] _1115;
    wire [7:0] _1110;
    wire [31:0] _1108;
    wire [23:0] _1109;
    wire [31:0] _1111;
    wire [31:0] _1112;
    wire [31:0] _1113;
    wire [24:0] _1114;
    wire [31:0] _1116;
    wire [63:0] _1105;
    wire [11:0] _1102;
    wire [15:0] _1097;
    wire [31:0] _1094;
    wire [31:0] _1095;
    wire [15:0] _1096;
    wire [31:0] _1098;
    wire [31:0] _1093;
    wire [31:0] _1099;
    wire [31:0] _1100;
    wire [19:0] _1101;
    wire [31:0] _1103;
    wire [31:0] _1091;
    wire [31:0] _1090;
    wire [31:0] _1092;
    wire [31:0] _1104;
    wire [383:0] _1087;
    wire [351:0] _1084;
    wire [191:0] _1081;
    wire [6:0] _1079;
    wire [7:0] _1074;
    wire [31:0] _1072;
    wire [23:0] _1073;
    wire [31:0] _1075;
    wire [31:0] _1076;
    wire [31:0] _1077;
    wire [24:0] _1078;
    wire [31:0] _1080;
    wire [31:0] _1069;
    wire [11:0] _1066;
    wire [15:0] _1061;
    wire [31:0] _1058;
    wire [31:0] _1059;
    wire [15:0] _1060;
    wire [31:0] _1062;
    wire [31:0] _1057;
    wire [31:0] _1063;
    wire [31:0] _1064;
    wire [19:0] _1065;
    wire [31:0] _1067;
    wire [31:0] _1055;
    wire [31:0] _1054;
    wire [31:0] _1056;
    wire [31:0] _1068;
    wire [319:0] _1049;
    wire [159:0] _1046;
    wire [6:0] _1044;
    wire [31:0] _1041;
    wire [31:0] _1042;
    wire [24:0] _1043;
    wire [31:0] _1045;
    wire [479:0] _1038;
    wire [511:0] _1039;
    wire [319:0] _1040;
    wire [511:0] _1047;
    wire [159:0] _1048;
    wire [511:0] _1050;
    wire [479:0] _1051;
    wire [7:0] _1036;
    wire [11:0] _1031;
    wire [31:0] _1027;
    wire [31:0] _1028;
    wire [31:0] _1029;
    wire [19:0] _1030;
    wire [31:0] _1032;
    wire [31:0] _1033;
    wire [15:0] _1025;
    wire [31:0] _1021;
    wire [31:0] _1020;
    wire [31:0] _1022;
    wire [351:0] _1015;
    wire [223:0] _1012;
    wire [6:0] _1010;
    wire [31:0] _1007;
    wire [31:0] _1008;
    wire [24:0] _1009;
    wire [31:0] _1011;
    wire [95:0] _1004;
    wire [383:0] _1003;
    wire [511:0] _1005;
    wire [255:0] _1006;
    wire [511:0] _1013;
    wire [127:0] _1014;
    wire [511:0] _1016;
    wire [479:0] _1017;
    wire [7:0] _1001;
    wire [11:0] _996;
    wire [31:0] _992;
    wire [31:0] _993;
    wire [31:0] _994;
    wire [19:0] _995;
    wire [31:0] _997;
    wire [31:0] _998;
    wire [15:0] _990;
    wire [31:0] _986;
    wire [31:0] _985;
    wire [31:0] _987;
    wire [447:0] _982;
    wire [319:0] _979;
    wire [191:0] _976;
    wire [6:0] _974;
    wire [7:0] _969;
    wire [31:0] _967;
    wire [23:0] _968;
    wire [31:0] _970;
    wire [31:0] _971;
    wire [31:0] _972;
    wire [24:0] _973;
    wire [31:0] _975;
    wire [63:0] _964;
    wire [11:0] _961;
    wire [15:0] _956;
    wire [31:0] _953;
    wire [31:0] _954;
    wire [15:0] _955;
    wire [31:0] _957;
    wire [31:0] _952;
    wire [31:0] _958;
    wire [31:0] _959;
    wire [19:0] _960;
    wire [31:0] _962;
    wire [31:0] _950;
    wire [31:0] _949;
    wire [31:0] _951;
    wire [31:0] _963;
    wire [415:0] _946;
    wire [287:0] _943;
    wire [159:0] _940;
    wire [6:0] _938;
    wire [7:0] _933;
    wire [31:0] _931;
    wire [23:0] _932;
    wire [31:0] _934;
    wire [31:0] _935;
    wire [31:0] _936;
    wire [24:0] _937;
    wire [31:0] _939;
    wire [31:0] _928;
    wire [11:0] _925;
    wire [15:0] _920;
    wire [31:0] _917;
    wire [31:0] _918;
    wire [15:0] _919;
    wire [31:0] _921;
    wire [31:0] _916;
    wire [31:0] _922;
    wire [31:0] _923;
    wire [19:0] _924;
    wire [31:0] _926;
    wire [31:0] _914;
    wire [31:0] _913;
    wire [31:0] _915;
    wire [31:0] _927;
    wire [383:0] _910;
    wire [255:0] _907;
    wire [127:0] _904;
    wire [6:0] _902;
    wire [7:0] _897;
    wire [31:0] _895;
    wire [23:0] _896;
    wire [31:0] _898;
    wire [31:0] _899;
    wire [31:0] _900;
    wire [24:0] _901;
    wire [31:0] _903;
    wire [11:0] _890;
    wire [15:0] _885;
    wire [31:0] _882;
    wire [31:0] _883;
    wire [15:0] _884;
    wire [31:0] _886;
    wire [31:0] _881;
    wire [31:0] _887;
    wire [31:0] _888;
    wire [19:0] _889;
    wire [31:0] _891;
    wire [31:0] _879;
    wire [31:0] _878;
    wire [31:0] _880;
    wire [31:0] _892;
    wire [447:0] _875;
    wire [287:0] _872;
    wire [127:0] _869;
    wire [6:0] _867;
    wire [7:0] _862;
    wire [31:0] _860;
    wire [23:0] _861;
    wire [31:0] _863;
    wire [31:0] _864;
    wire [31:0] _865;
    wire [24:0] _866;
    wire [31:0] _868;
    wire [95:0] _857;
    wire [11:0] _854;
    wire [15:0] _849;
    wire [31:0] _846;
    wire [31:0] _847;
    wire [15:0] _848;
    wire [31:0] _850;
    wire [31:0] _845;
    wire [31:0] _851;
    wire [31:0] _852;
    wire [19:0] _853;
    wire [31:0] _855;
    wire [31:0] _843;
    wire [31:0] _842;
    wire [31:0] _844;
    wire [31:0] _856;
    wire [415:0] _839;
    wire [255:0] _836;
    wire [223:0] _833;
    wire [6:0] _831;
    wire [7:0] _826;
    wire [31:0] _824;
    wire [23:0] _825;
    wire [31:0] _827;
    wire [31:0] _828;
    wire [31:0] _829;
    wire [24:0] _830;
    wire [31:0] _832;
    wire [63:0] _821;
    wire [11:0] _818;
    wire [15:0] _813;
    wire [31:0] _810;
    wire [31:0] _811;
    wire [15:0] _812;
    wire [31:0] _814;
    wire [31:0] _809;
    wire [31:0] _815;
    wire [31:0] _816;
    wire [19:0] _817;
    wire [31:0] _819;
    wire [31:0] _807;
    wire [31:0] _806;
    wire [31:0] _808;
    wire [31:0] _820;
    wire [383:0] _803;
    wire [351:0] _800;
    wire [191:0] _797;
    wire [6:0] _795;
    wire [7:0] _790;
    wire [31:0] _788;
    wire [23:0] _789;
    wire [31:0] _791;
    wire [31:0] _792;
    wire [31:0] _793;
    wire [24:0] _794;
    wire [31:0] _796;
    wire [31:0] _785;
    wire [11:0] _782;
    wire [15:0] _777;
    wire [31:0] _774;
    wire [31:0] _775;
    wire [15:0] _776;
    wire [31:0] _778;
    wire [31:0] _773;
    wire [31:0] _779;
    wire [31:0] _780;
    wire [19:0] _781;
    wire [31:0] _783;
    wire [31:0] _771;
    wire [31:0] _770;
    wire [31:0] _772;
    wire [31:0] _784;
    wire [319:0] _765;
    wire [159:0] _762;
    wire [6:0] _760;
    wire [31:0] _757;
    wire [31:0] _758;
    wire [24:0] _759;
    wire [31:0] _761;
    wire [479:0] _754;
    wire [511:0] _755;
    wire [319:0] _756;
    wire [511:0] _763;
    wire [159:0] _764;
    wire [511:0] _766;
    wire [479:0] _767;
    wire [7:0] _752;
    wire [11:0] _747;
    wire [31:0] _743;
    wire [31:0] _744;
    wire [31:0] _745;
    wire [19:0] _746;
    wire [31:0] _748;
    wire [31:0] _749;
    wire [15:0] _741;
    wire [31:0] _737;
    wire [31:0] _736;
    wire [31:0] _738;
    wire [351:0] _731;
    wire [223:0] _728;
    wire [6:0] _726;
    wire [31:0] _723;
    wire [31:0] _724;
    wire [24:0] _725;
    wire [31:0] _727;
    wire [95:0] _720;
    wire [383:0] _719;
    wire [511:0] _721;
    wire [255:0] _722;
    wire [511:0] _729;
    wire [127:0] _730;
    wire [511:0] _732;
    wire [479:0] _733;
    wire [7:0] _717;
    wire [11:0] _712;
    wire [31:0] _708;
    wire [31:0] _709;
    wire [31:0] _710;
    wire [19:0] _711;
    wire [31:0] _713;
    wire [31:0] _714;
    wire [15:0] _706;
    wire [31:0] _702;
    wire [31:0] _701;
    wire [31:0] _703;
    wire [447:0] _698;
    wire [319:0] _695;
    wire [191:0] _692;
    wire [6:0] _690;
    wire [7:0] _685;
    wire [31:0] _683;
    wire [23:0] _684;
    wire [31:0] _686;
    wire [31:0] _687;
    wire [31:0] _688;
    wire [24:0] _689;
    wire [31:0] _691;
    wire [63:0] _680;
    wire [11:0] _677;
    wire [15:0] _672;
    wire [31:0] _669;
    wire [31:0] _670;
    wire [15:0] _671;
    wire [31:0] _673;
    wire [31:0] _668;
    wire [31:0] _674;
    wire [31:0] _675;
    wire [19:0] _676;
    wire [31:0] _678;
    wire [31:0] _666;
    wire [31:0] _665;
    wire [31:0] _667;
    wire [31:0] _679;
    wire [415:0] _662;
    wire [287:0] _659;
    wire [159:0] _656;
    wire [6:0] _654;
    wire [7:0] _649;
    wire [31:0] _647;
    wire [23:0] _648;
    wire [31:0] _650;
    wire [31:0] _651;
    wire [31:0] _652;
    wire [24:0] _653;
    wire [31:0] _655;
    wire [31:0] _644;
    wire [11:0] _641;
    wire [15:0] _636;
    wire [31:0] _633;
    wire [31:0] _634;
    wire [15:0] _635;
    wire [31:0] _637;
    wire [31:0] _632;
    wire [31:0] _638;
    wire [31:0] _639;
    wire [19:0] _640;
    wire [31:0] _642;
    wire [31:0] _630;
    wire [31:0] _629;
    wire [31:0] _631;
    wire [31:0] _643;
    wire [383:0] _626;
    wire [255:0] _623;
    wire [127:0] _620;
    wire [6:0] _618;
    wire [7:0] _613;
    wire [31:0] _611;
    wire [23:0] _612;
    wire [31:0] _614;
    wire [31:0] _615;
    wire [31:0] _616;
    wire [24:0] _617;
    wire [31:0] _619;
    wire [11:0] _606;
    wire [15:0] _601;
    wire [31:0] _598;
    wire [31:0] _599;
    wire [15:0] _600;
    wire [31:0] _602;
    wire [31:0] _597;
    wire [31:0] _603;
    wire [31:0] _604;
    wire [19:0] _605;
    wire [31:0] _607;
    wire [31:0] _595;
    wire [31:0] _594;
    wire [31:0] _596;
    wire [31:0] _608;
    wire [447:0] _591;
    wire [287:0] _588;
    wire [127:0] _585;
    wire [6:0] _583;
    wire [7:0] _578;
    wire [31:0] _576;
    wire [23:0] _577;
    wire [31:0] _579;
    wire [31:0] _580;
    wire [31:0] _581;
    wire [24:0] _582;
    wire [31:0] _584;
    wire [95:0] _573;
    wire [11:0] _570;
    wire [15:0] _565;
    wire [31:0] _562;
    wire [31:0] _563;
    wire [15:0] _564;
    wire [31:0] _566;
    wire [31:0] _561;
    wire [31:0] _567;
    wire [31:0] _568;
    wire [19:0] _569;
    wire [31:0] _571;
    wire [31:0] _559;
    wire [31:0] _558;
    wire [31:0] _560;
    wire [31:0] _572;
    wire [415:0] _555;
    wire [255:0] _552;
    wire [223:0] _549;
    wire [6:0] _547;
    wire [7:0] _542;
    wire [31:0] _540;
    wire [23:0] _541;
    wire [31:0] _543;
    wire [31:0] _544;
    wire [31:0] _545;
    wire [24:0] _546;
    wire [31:0] _548;
    wire [63:0] _537;
    wire [11:0] _534;
    wire [15:0] _529;
    wire [31:0] _526;
    wire [31:0] _527;
    wire [15:0] _528;
    wire [31:0] _530;
    wire [31:0] _525;
    wire [31:0] _531;
    wire [31:0] _532;
    wire [19:0] _533;
    wire [31:0] _535;
    wire [31:0] _523;
    wire [31:0] _522;
    wire [31:0] _524;
    wire [31:0] _536;
    wire [383:0] _519;
    wire [351:0] _516;
    wire [191:0] _513;
    wire [6:0] _511;
    wire [7:0] _506;
    wire [31:0] _504;
    wire [23:0] _505;
    wire [31:0] _507;
    wire [31:0] _508;
    wire [31:0] _509;
    wire [24:0] _510;
    wire [31:0] _512;
    wire [31:0] _501;
    wire [11:0] _498;
    wire [15:0] _493;
    wire [31:0] _490;
    wire [31:0] _491;
    wire [15:0] _492;
    wire [31:0] _494;
    wire [31:0] _489;
    wire [31:0] _495;
    wire [31:0] _496;
    wire [19:0] _497;
    wire [31:0] _499;
    wire [31:0] _487;
    wire [31:0] _486;
    wire [31:0] _488;
    wire [31:0] _500;
    wire [319:0] _481;
    wire [159:0] _478;
    wire [6:0] _476;
    wire [31:0] _473;
    wire [31:0] _474;
    wire [24:0] _475;
    wire [31:0] _477;
    wire [479:0] _470;
    wire [511:0] _471;
    wire [319:0] _472;
    wire [511:0] _479;
    wire [159:0] _480;
    wire [511:0] _482;
    wire [479:0] _483;
    wire [7:0] _468;
    wire [11:0] _463;
    wire [31:0] _459;
    wire [31:0] _460;
    wire [31:0] _461;
    wire [19:0] _462;
    wire [31:0] _464;
    wire [31:0] _465;
    wire [15:0] _457;
    wire [31:0] _453;
    wire [31:0] _452;
    wire [31:0] _454;
    wire [351:0] _447;
    wire [223:0] _444;
    wire [6:0] _442;
    wire [31:0] _439;
    wire [31:0] _440;
    wire [24:0] _441;
    wire [31:0] _443;
    wire [95:0] _436;
    wire [383:0] _435;
    wire [511:0] _437;
    wire [255:0] _438;
    wire [511:0] _445;
    wire [127:0] _446;
    wire [511:0] _448;
    wire [479:0] _449;
    wire [7:0] _433;
    wire [11:0] _428;
    wire [31:0] _424;
    wire [31:0] _425;
    wire [31:0] _426;
    wire [19:0] _427;
    wire [31:0] _429;
    wire [31:0] _430;
    wire [15:0] _422;
    wire [31:0] _418;
    wire [31:0] _417;
    wire [31:0] _419;
    wire [447:0] _414;
    wire [319:0] _411;
    wire [191:0] _408;
    wire [6:0] _406;
    wire [7:0] _401;
    wire [31:0] _399;
    wire [23:0] _400;
    wire [31:0] _402;
    wire [31:0] _403;
    wire [31:0] _404;
    wire [24:0] _405;
    wire [31:0] _407;
    wire [63:0] _396;
    wire [11:0] _393;
    wire [15:0] _388;
    wire [31:0] _385;
    wire [31:0] _386;
    wire [15:0] _387;
    wire [31:0] _389;
    wire [31:0] _384;
    wire [31:0] _390;
    wire [31:0] _391;
    wire [19:0] _392;
    wire [31:0] _394;
    wire [31:0] _382;
    wire [31:0] _381;
    wire [31:0] _383;
    wire [31:0] _395;
    wire [415:0] _378;
    wire [287:0] _375;
    wire [159:0] _372;
    wire [6:0] _370;
    wire [7:0] _365;
    wire [31:0] _363;
    wire [23:0] _364;
    wire [31:0] _366;
    wire [31:0] _367;
    wire [31:0] _368;
    wire [24:0] _369;
    wire [31:0] _371;
    wire [31:0] _360;
    wire [11:0] _357;
    wire [15:0] _352;
    wire [31:0] _349;
    wire [31:0] _350;
    wire [15:0] _351;
    wire [31:0] _353;
    wire [31:0] _348;
    wire [31:0] _354;
    wire [31:0] _355;
    wire [19:0] _356;
    wire [31:0] _358;
    wire [31:0] _346;
    wire [31:0] _345;
    wire [31:0] _347;
    wire [31:0] _359;
    wire [383:0] _342;
    wire [255:0] _339;
    wire [127:0] _336;
    wire [6:0] _334;
    wire [7:0] _329;
    wire [31:0] _327;
    wire [23:0] _328;
    wire [31:0] _330;
    wire [31:0] _331;
    wire [31:0] _332;
    wire [24:0] _333;
    wire [31:0] _335;
    wire [11:0] _322;
    wire [15:0] _317;
    wire [31:0] _314;
    wire [31:0] _315;
    wire [15:0] _316;
    wire [31:0] _318;
    wire [31:0] _313;
    wire [31:0] _319;
    wire [31:0] _320;
    wire [19:0] _321;
    wire [31:0] _323;
    wire [31:0] _311;
    wire [31:0] _310;
    wire [31:0] _312;
    wire [31:0] _324;
    wire [447:0] _307;
    wire [287:0] _304;
    wire [127:0] _301;
    wire [6:0] _299;
    wire [7:0] _294;
    wire [31:0] _292;
    wire [23:0] _293;
    wire [31:0] _295;
    wire [31:0] _296;
    wire [31:0] _297;
    wire [24:0] _298;
    wire [31:0] _300;
    wire [95:0] _289;
    wire [11:0] _286;
    wire [15:0] _281;
    wire [31:0] _278;
    wire [31:0] _279;
    wire [15:0] _280;
    wire [31:0] _282;
    wire [31:0] _277;
    wire [31:0] _283;
    wire [31:0] _284;
    wire [19:0] _285;
    wire [31:0] _287;
    wire [31:0] _275;
    wire [31:0] _274;
    wire [31:0] _276;
    wire [31:0] _288;
    wire [415:0] _271;
    wire [255:0] _268;
    wire [223:0] _265;
    wire [6:0] _263;
    wire [7:0] _258;
    wire [31:0] _256;
    wire [23:0] _257;
    wire [31:0] _259;
    wire [31:0] _260;
    wire [31:0] _261;
    wire [24:0] _262;
    wire [31:0] _264;
    wire [63:0] _253;
    wire [11:0] _250;
    wire [15:0] _245;
    wire [31:0] _242;
    wire [31:0] _243;
    wire [15:0] _244;
    wire [31:0] _246;
    wire [31:0] _241;
    wire [31:0] _247;
    wire [31:0] _248;
    wire [19:0] _249;
    wire [31:0] _251;
    wire [31:0] _239;
    wire [31:0] _238;
    wire [31:0] _240;
    wire [31:0] _252;
    wire [383:0] _235;
    wire [351:0] _232;
    wire [191:0] _229;
    wire [6:0] _227;
    wire [7:0] _222;
    wire [31:0] _220;
    wire [23:0] _221;
    wire [31:0] _223;
    wire [31:0] _224;
    wire [31:0] _225;
    wire [24:0] _226;
    wire [31:0] _228;
    wire [31:0] _217;
    wire [11:0] _214;
    wire [15:0] _209;
    wire [31:0] _206;
    wire [31:0] _207;
    wire [15:0] _208;
    wire [31:0] _210;
    wire [31:0] _205;
    wire [31:0] _211;
    wire [31:0] _212;
    wire [19:0] _213;
    wire [31:0] _215;
    wire [31:0] _203;
    wire [31:0] _202;
    wire [31:0] _204;
    wire [31:0] _216;
    wire [319:0] _197;
    wire [159:0] _194;
    wire [6:0] _192;
    wire [31:0] _189;
    wire [31:0] _190;
    wire [24:0] _191;
    wire [31:0] _193;
    wire [479:0] _186;
    wire [511:0] _187;
    wire [319:0] _188;
    wire [511:0] _195;
    wire [159:0] _196;
    wire [511:0] _198;
    wire [479:0] _199;
    wire [7:0] _184;
    wire [11:0] _179;
    wire [31:0] _175;
    wire [31:0] _176;
    wire [31:0] _177;
    wire [19:0] _178;
    wire [31:0] _180;
    wire [31:0] _181;
    wire [15:0] _173;
    wire [31:0] _169;
    wire [31:0] _168;
    wire [31:0] _170;
    wire [351:0] _163;
    wire [223:0] _160;
    wire [6:0] _158;
    wire [31:0] _155;
    wire [31:0] _156;
    wire [24:0] _157;
    wire [31:0] _159;
    wire [95:0] _152;
    wire [383:0] _151;
    wire [511:0] _153;
    wire [255:0] _154;
    wire [511:0] _161;
    wire [127:0] _162;
    wire [511:0] _164;
    wire [479:0] _165;
    wire [7:0] _149;
    wire [11:0] _144;
    wire [31:0] _140;
    wire [31:0] _141;
    wire [31:0] _142;
    wire [19:0] _143;
    wire [31:0] _145;
    wire [31:0] _146;
    wire [15:0] _138;
    wire [31:0] _134;
    wire [31:0] _133;
    wire [31:0] _135;
    wire [447:0] _130;
    wire [319:0] _127;
    wire [191:0] _124;
    wire [6:0] _122;
    wire [7:0] _117;
    wire [31:0] _115;
    wire [23:0] _116;
    wire [31:0] _118;
    wire [31:0] _119;
    wire [31:0] _120;
    wire [24:0] _121;
    wire [31:0] _123;
    wire [63:0] _112;
    wire [11:0] _109;
    wire [15:0] _104;
    wire [31:0] _101;
    wire [31:0] _102;
    wire [15:0] _103;
    wire [31:0] _105;
    wire [31:0] _100;
    wire [31:0] _106;
    wire [31:0] _107;
    wire [19:0] _108;
    wire [31:0] _110;
    wire [31:0] _98;
    wire [31:0] _97;
    wire [31:0] _99;
    wire [31:0] _111;
    wire [415:0] _94;
    wire [287:0] _91;
    wire [159:0] _88;
    wire [6:0] _86;
    wire [7:0] _81;
    wire [31:0] _79;
    wire [23:0] _80;
    wire [31:0] _82;
    wire [31:0] _83;
    wire [31:0] _84;
    wire [24:0] _85;
    wire [31:0] _87;
    wire [31:0] _76;
    wire [11:0] _73;
    wire [15:0] _68;
    wire [31:0] _65;
    wire [31:0] _66;
    wire [15:0] _67;
    wire [31:0] _69;
    wire [31:0] _64;
    wire [31:0] _70;
    wire [31:0] _71;
    wire [19:0] _72;
    wire [31:0] _74;
    wire [31:0] _62;
    wire [31:0] _61;
    wire [31:0] _63;
    wire [31:0] _75;
    wire [383:0] _58;
    wire [255:0] _55;
    wire [127:0] _52;
    wire [6:0] _50;
    wire [7:0] _45;
    wire [31:0] _43;
    wire [23:0] _44;
    wire [31:0] _46;
    wire [31:0] _47;
    wire [31:0] _48;
    wire [24:0] _49;
    wire [31:0] _51;
    wire [11:0] _38;
    wire [15:0] _33;
    wire [31:0] _30;
    wire [31:0] _31;
    wire [15:0] _32;
    wire [31:0] _34;
    wire [31:0] _29;
    wire [31:0] _35;
    wire [31:0] _36;
    wire [19:0] _37;
    wire [31:0] _39;
    wire [31:0] _27;
    wire [31:0] _26;
    wire [31:0] _28;
    wire [31:0] _40;
    wire [479:0] _25;
    wire [511:0] _41;
    wire [351:0] _42;
    wire [511:0] _53;
    wire [223:0] _54;
    wire [511:0] _56;
    wire [95:0] _57;
    wire [511:0] _59;
    wire [447:0] _60;
    wire [511:0] _77;
    wire [319:0] _78;
    wire [511:0] _89;
    wire [191:0] _90;
    wire [511:0] _92;
    wire [63:0] _93;
    wire [511:0] _95;
    wire [415:0] _96;
    wire [511:0] _113;
    wire [287:0] _114;
    wire [511:0] _125;
    wire [159:0] _126;
    wire [511:0] _128;
    wire [31:0] _129;
    wire [511:0] _131;
    wire [31:0] _132;
    wire [31:0] _136;
    wire [15:0] _137;
    wire [31:0] _139;
    wire [31:0] _147;
    wire [23:0] _148;
    wire [31:0] _150;
    wire [511:0] _166;
    wire [31:0] _167;
    wire [31:0] _171;
    wire [15:0] _172;
    wire [31:0] _174;
    wire [31:0] _182;
    wire [23:0] _183;
    wire [31:0] _185;
    wire [511:0] _200;
    wire [447:0] _201;
    wire [511:0] _218;
    wire [287:0] _219;
    wire [511:0] _230;
    wire [127:0] _231;
    wire [511:0] _233;
    wire [95:0] _234;
    wire [511:0] _236;
    wire [415:0] _237;
    wire [511:0] _254;
    wire [255:0] _255;
    wire [511:0] _266;
    wire [223:0] _267;
    wire [511:0] _269;
    wire [63:0] _270;
    wire [511:0] _272;
    wire [383:0] _273;
    wire [511:0] _290;
    wire [351:0] _291;
    wire [511:0] _302;
    wire [191:0] _303;
    wire [511:0] _305;
    wire [31:0] _306;
    wire [511:0] _308;
    wire [479:0] _309;
    wire [511:0] _325;
    wire [351:0] _326;
    wire [511:0] _337;
    wire [223:0] _338;
    wire [511:0] _340;
    wire [95:0] _341;
    wire [511:0] _343;
    wire [447:0] _344;
    wire [511:0] _361;
    wire [319:0] _362;
    wire [511:0] _373;
    wire [191:0] _374;
    wire [511:0] _376;
    wire [63:0] _377;
    wire [511:0] _379;
    wire [415:0] _380;
    wire [511:0] _397;
    wire [287:0] _398;
    wire [511:0] _409;
    wire [159:0] _410;
    wire [511:0] _412;
    wire [31:0] _413;
    wire [511:0] _415;
    wire [31:0] _416;
    wire [31:0] _420;
    wire [15:0] _421;
    wire [31:0] _423;
    wire [31:0] _431;
    wire [23:0] _432;
    wire [31:0] _434;
    wire [511:0] _450;
    wire [31:0] _451;
    wire [31:0] _455;
    wire [15:0] _456;
    wire [31:0] _458;
    wire [31:0] _466;
    wire [23:0] _467;
    wire [31:0] _469;
    wire [511:0] _484;
    wire [447:0] _485;
    wire [511:0] _502;
    wire [287:0] _503;
    wire [511:0] _514;
    wire [127:0] _515;
    wire [511:0] _517;
    wire [95:0] _518;
    wire [511:0] _520;
    wire [415:0] _521;
    wire [511:0] _538;
    wire [255:0] _539;
    wire [511:0] _550;
    wire [223:0] _551;
    wire [511:0] _553;
    wire [63:0] _554;
    wire [511:0] _556;
    wire [383:0] _557;
    wire [511:0] _574;
    wire [351:0] _575;
    wire [511:0] _586;
    wire [191:0] _587;
    wire [511:0] _589;
    wire [31:0] _590;
    wire [511:0] _592;
    wire [479:0] _593;
    wire [511:0] _609;
    wire [351:0] _610;
    wire [511:0] _621;
    wire [223:0] _622;
    wire [511:0] _624;
    wire [95:0] _625;
    wire [511:0] _627;
    wire [447:0] _628;
    wire [511:0] _645;
    wire [319:0] _646;
    wire [511:0] _657;
    wire [191:0] _658;
    wire [511:0] _660;
    wire [63:0] _661;
    wire [511:0] _663;
    wire [415:0] _664;
    wire [511:0] _681;
    wire [287:0] _682;
    wire [511:0] _693;
    wire [159:0] _694;
    wire [511:0] _696;
    wire [31:0] _697;
    wire [511:0] _699;
    wire [31:0] _700;
    wire [31:0] _704;
    wire [15:0] _705;
    wire [31:0] _707;
    wire [31:0] _715;
    wire [23:0] _716;
    wire [31:0] _718;
    wire [511:0] _734;
    wire [31:0] _735;
    wire [31:0] _739;
    wire [15:0] _740;
    wire [31:0] _742;
    wire [31:0] _750;
    wire [23:0] _751;
    wire [31:0] _753;
    wire [511:0] _768;
    wire [447:0] _769;
    wire [511:0] _786;
    wire [287:0] _787;
    wire [511:0] _798;
    wire [127:0] _799;
    wire [511:0] _801;
    wire [95:0] _802;
    wire [511:0] _804;
    wire [415:0] _805;
    wire [511:0] _822;
    wire [255:0] _823;
    wire [511:0] _834;
    wire [223:0] _835;
    wire [511:0] _837;
    wire [63:0] _838;
    wire [511:0] _840;
    wire [383:0] _841;
    wire [511:0] _858;
    wire [351:0] _859;
    wire [511:0] _870;
    wire [191:0] _871;
    wire [511:0] _873;
    wire [31:0] _874;
    wire [511:0] _876;
    wire [479:0] _877;
    wire [511:0] _893;
    wire [351:0] _894;
    wire [511:0] _905;
    wire [223:0] _906;
    wire [511:0] _908;
    wire [95:0] _909;
    wire [511:0] _911;
    wire [447:0] _912;
    wire [511:0] _929;
    wire [319:0] _930;
    wire [511:0] _941;
    wire [191:0] _942;
    wire [511:0] _944;
    wire [63:0] _945;
    wire [511:0] _947;
    wire [415:0] _948;
    wire [511:0] _965;
    wire [287:0] _966;
    wire [511:0] _977;
    wire [159:0] _978;
    wire [511:0] _980;
    wire [31:0] _981;
    wire [511:0] _983;
    wire [31:0] _984;
    wire [31:0] _988;
    wire [15:0] _989;
    wire [31:0] _991;
    wire [31:0] _999;
    wire [23:0] _1000;
    wire [31:0] _1002;
    wire [511:0] _1018;
    wire [31:0] _1019;
    wire [31:0] _1023;
    wire [15:0] _1024;
    wire [31:0] _1026;
    wire [31:0] _1034;
    wire [23:0] _1035;
    wire [31:0] _1037;
    wire [511:0] _1052;
    wire [447:0] _1053;
    wire [511:0] _1070;
    wire [287:0] _1071;
    wire [511:0] _1082;
    wire [127:0] _1083;
    wire [511:0] _1085;
    wire [95:0] _1086;
    wire [511:0] _1088;
    wire [415:0] _1089;
    wire [511:0] _1106;
    wire [255:0] _1107;
    wire [511:0] _1118;
    wire [223:0] _1119;
    wire [511:0] _1121;
    wire [63:0] _1122;
    wire [511:0] _1124;
    wire [383:0] _1125;
    wire [511:0] _1142;
    wire [351:0] _1143;
    wire [511:0] _1154;
    wire [191:0] _1155;
    wire [511:0] _1157;
    wire [31:0] _1158;
    wire [511:0] _1160;
    wire [479:0] _1161;
    wire [511:0] _1177;
    wire [351:0] _1178;
    wire [511:0] _1189;
    wire [223:0] _1190;
    wire [511:0] _1192;
    wire [95:0] _1193;
    wire [511:0] _1195;
    wire [447:0] _1196;
    wire [511:0] _1213;
    wire [319:0] _1214;
    wire [511:0] _1225;
    wire [191:0] _1226;
    wire [511:0] _1228;
    wire [63:0] _1229;
    wire [511:0] _1231;
    wire [415:0] _1232;
    wire [511:0] _1249;
    wire [287:0] _1250;
    wire [511:0] _1261;
    wire [159:0] _1262;
    wire [511:0] _1264;
    wire [31:0] _1265;
    wire [511:0] _1267;
    wire [31:0] _1268;
    wire [31:0] _1272;
    wire [15:0] _1273;
    wire [31:0] _1275;
    wire [31:0] _1283;
    wire [23:0] _1284;
    wire [31:0] _1286;
    wire [511:0] _1302;
    wire [31:0] _1303;
    wire [31:0] _1307;
    wire [15:0] _1308;
    wire [31:0] _1310;
    wire [31:0] _1318;
    wire [23:0] _1319;
    wire [31:0] _1321;
    wire [511:0] _1336;
    wire [447:0] _1337;
    wire [511:0] _1354;
    wire [287:0] _1355;
    wire [511:0] _1366;
    wire [127:0] _1367;
    wire [511:0] _1369;
    wire [95:0] _1370;
    wire [511:0] _1372;
    wire [415:0] _1373;
    wire [511:0] _1390;
    wire [255:0] _1391;
    wire [511:0] _1402;
    wire [223:0] _1403;
    wire [511:0] _1405;
    wire [63:0] _1406;
    wire [511:0] _1408;
    wire [383:0] _1409;
    wire [511:0] _1426;
    wire [351:0] _1427;
    wire [511:0] _1438;
    wire [191:0] _1439;
    wire [511:0] _1441;
    wire [31:0] _1442;
    wire [511:0] _1444;
    wire [479:0] _1445;
    wire [511:0] _1461;
    wire [351:0] _1462;
    wire [511:0] _1473;
    wire [223:0] _1474;
    wire [511:0] _1476;
    wire [95:0] _1477;
    wire [511:0] _1479;
    wire [447:0] _1480;
    wire [511:0] _1497;
    wire [319:0] _1498;
    wire [511:0] _1509;
    wire [191:0] _1510;
    wire [511:0] _1512;
    wire [63:0] _1513;
    wire [511:0] _1515;
    wire [415:0] _1516;
    wire [511:0] _1533;
    wire [287:0] _1534;
    wire [511:0] _1545;
    wire [159:0] _1546;
    wire [511:0] _1548;
    wire [31:0] _1549;
    wire [511:0] _1551;
    wire [31:0] _1552;
    wire [31:0] _1556;
    wire [15:0] _1557;
    wire [31:0] _1559;
    wire [31:0] _1567;
    wire [23:0] _1568;
    wire [31:0] _1570;
    wire [511:0] _1586;
    wire [31:0] _1587;
    wire [31:0] _1591;
    wire [15:0] _1592;
    wire [31:0] _1594;
    wire [31:0] _1602;
    wire [23:0] _1603;
    wire [31:0] _1605;
    wire [511:0] _1620;
    wire [447:0] _1621;
    wire [511:0] _1638;
    wire [287:0] _1639;
    wire [511:0] _1650;
    wire [127:0] _1651;
    wire [511:0] _1653;
    wire [95:0] _1654;
    wire [511:0] _1656;
    wire [415:0] _1657;
    wire [511:0] _1674;
    wire [255:0] _1675;
    wire [511:0] _1686;
    wire [223:0] _1687;
    wire [511:0] _1689;
    wire [63:0] _1690;
    wire [511:0] _1692;
    wire [383:0] _1693;
    wire [511:0] _1710;
    wire [351:0] _1711;
    wire [511:0] _1722;
    wire [191:0] _1723;
    wire [511:0] _1725;
    wire [31:0] _1726;
    wire [511:0] _1728;
    wire [479:0] _1729;
    wire [511:0] _1745;
    wire [351:0] _1746;
    wire [511:0] _1757;
    wire [223:0] _1758;
    wire [511:0] _1760;
    wire [95:0] _1761;
    wire [511:0] _1763;
    wire [447:0] _1764;
    wire [511:0] _1781;
    wire [319:0] _1782;
    wire [511:0] _1793;
    wire [191:0] _1794;
    wire [511:0] _1796;
    wire [63:0] _1797;
    wire [511:0] _1799;
    wire [415:0] _1800;
    wire [511:0] _1817;
    wire [287:0] _1818;
    wire [511:0] _1829;
    wire [159:0] _1830;
    wire [511:0] _1832;
    wire [31:0] _1833;
    wire [511:0] _1835;
    wire [31:0] _1836;
    wire [31:0] _1840;
    wire [15:0] _1841;
    wire [31:0] _1843;
    wire [31:0] _1851;
    wire [23:0] _1852;
    wire [31:0] _1854;
    wire [511:0] _1870;
    wire [31:0] _1871;
    wire [31:0] _1875;
    wire [15:0] _1876;
    wire [31:0] _1878;
    wire [31:0] _1886;
    wire [23:0] _1887;
    wire [31:0] _1889;
    wire [511:0] _1904;
    wire [447:0] _1905;
    wire [511:0] _1922;
    wire [287:0] _1923;
    wire [511:0] _1934;
    wire [127:0] _1935;
    wire [511:0] _1937;
    wire [95:0] _1938;
    wire [511:0] _1940;
    wire [415:0] _1941;
    wire [511:0] _1958;
    wire [255:0] _1959;
    wire [511:0] _1970;
    wire [223:0] _1971;
    wire [511:0] _1973;
    wire [63:0] _1974;
    wire [511:0] _1976;
    wire [383:0] _1977;
    wire [511:0] _1994;
    wire [351:0] _1995;
    wire [511:0] _2006;
    wire [191:0] _2007;
    wire [511:0] _2009;
    wire [31:0] _2010;
    wire [511:0] _2012;
    wire [479:0] _2013;
    wire [511:0] _2029;
    wire [351:0] _2030;
    wire [511:0] _2041;
    wire [223:0] _2042;
    wire [511:0] _2044;
    wire [95:0] _2045;
    wire [511:0] _2047;
    wire [447:0] _2048;
    wire [511:0] _2065;
    wire [319:0] _2066;
    wire [511:0] _2077;
    wire [191:0] _2078;
    wire [511:0] _2080;
    wire [63:0] _2081;
    wire [511:0] _2083;
    wire [415:0] _2084;
    wire [511:0] _2101;
    wire [287:0] _2102;
    wire [511:0] _2113;
    wire [159:0] _2114;
    wire [511:0] _2116;
    wire [31:0] _2117;
    wire [511:0] _2119;
    wire [31:0] _2120;
    wire [31:0] _2124;
    wire [15:0] _2125;
    wire [31:0] _2127;
    wire [31:0] _2135;
    wire [23:0] _2136;
    wire [31:0] _2138;
    wire [511:0] _2154;
    wire [31:0] _2155;
    wire [31:0] _2159;
    wire [15:0] _2160;
    wire [31:0] _2162;
    wire [31:0] _2170;
    wire [23:0] _2171;
    wire [31:0] _2173;
    wire [511:0] _2188;
    wire [447:0] _2189;
    wire [511:0] _2206;
    wire [287:0] _2207;
    wire [511:0] _2218;
    wire [127:0] _2219;
    wire [511:0] _2221;
    wire [95:0] _2222;
    wire [511:0] _2224;
    wire [415:0] _2225;
    wire [511:0] _2242;
    wire [255:0] _2243;
    wire [511:0] _2254;
    wire [223:0] _2255;
    wire [511:0] _2257;
    wire [63:0] _2258;
    wire [511:0] _2260;
    wire [383:0] _2261;
    wire [511:0] _2278;
    wire [351:0] _2279;
    wire [511:0] _2290;
    wire [191:0] _2291;
    wire [511:0] _2293;
    wire [31:0] _2294;
    wire [511:0] _2296;
    wire [479:0] _2297;
    wire [511:0] _2313;
    wire [351:0] _2314;
    wire [511:0] _2325;
    wire [223:0] _2326;
    wire [511:0] _2328;
    wire [95:0] _2329;
    wire [511:0] _2331;
    wire [447:0] _2332;
    wire [511:0] _2349;
    wire [319:0] _2350;
    wire [511:0] _2361;
    wire [191:0] _2362;
    wire [511:0] _2364;
    wire [63:0] _2365;
    wire [511:0] _2367;
    wire [415:0] _2368;
    wire [511:0] _2385;
    wire [287:0] _2386;
    wire [511:0] _2397;
    wire [159:0] _2398;
    wire [511:0] _2400;
    wire [31:0] _2401;
    wire [511:0] _2403;
    wire [31:0] _2404;
    wire [31:0] _2408;
    wire [15:0] _2409;
    wire [31:0] _2411;
    wire [31:0] _2419;
    wire [23:0] _2420;
    wire [31:0] _2422;
    wire [511:0] _2438;
    wire [31:0] _2439;
    wire [31:0] _2443;
    wire [15:0] _2444;
    wire [31:0] _2446;
    wire [31:0] _2454;
    wire [23:0] _2455;
    wire [31:0] _2457;
    wire [511:0] _2472;
    wire [447:0] _2473;
    wire [511:0] _2490;
    wire [287:0] _2491;
    wire [511:0] _2502;
    wire [127:0] _2503;
    wire [511:0] _2505;
    wire [95:0] _2506;
    wire [511:0] _2508;
    wire [415:0] _2509;
    wire [511:0] _2526;
    wire [255:0] _2527;
    wire [511:0] _2538;
    wire [223:0] _2539;
    wire [511:0] _2541;
    wire [63:0] _2542;
    wire [511:0] _2544;
    wire [383:0] _2545;
    wire [511:0] _2562;
    wire [351:0] _2563;
    wire [511:0] _2574;
    wire [191:0] _2575;
    wire [511:0] _2577;
    wire [31:0] _2578;
    wire [511:0] _2580;
    wire [479:0] _2581;
    wire [511:0] _2597;
    wire [351:0] _2598;
    wire [511:0] _2609;
    wire [223:0] _2610;
    wire [511:0] _2612;
    wire [95:0] _2613;
    wire [511:0] _2615;
    wire [447:0] _2616;
    wire [511:0] _2633;
    wire [319:0] _2634;
    wire [511:0] _2645;
    wire [191:0] _2646;
    wire [511:0] _2648;
    wire [63:0] _2649;
    wire [511:0] _2651;
    wire [415:0] _2652;
    wire [511:0] _2669;
    wire [287:0] _2670;
    wire [511:0] _2681;
    wire [159:0] _2682;
    wire [511:0] _2684;
    wire [31:0] _2685;
    wire [511:0] _2687;
    wire [31:0] _2688;
    wire [31:0] _2692;
    wire [15:0] _2693;
    wire [31:0] _2695;
    wire [31:0] _2703;
    wire [23:0] _2704;
    wire [31:0] _2706;
    wire [511:0] _2722;
    wire [31:0] _2723;
    wire [31:0] _2727;
    wire [15:0] _2728;
    wire [31:0] _2730;
    wire [31:0] _2738;
    wire [23:0] _2739;
    wire [31:0] _2741;
    wire [511:0] _2756;
    wire [447:0] _2757;
    wire [511:0] _2774;
    wire [287:0] _2775;
    wire [511:0] _2786;
    wire [127:0] _2787;
    wire [511:0] _2789;
    wire [95:0] _2790;
    wire [511:0] _2792;
    wire [415:0] _2793;
    wire [511:0] _2810;
    wire [255:0] _2811;
    wire [511:0] _2822;
    wire [223:0] _2823;
    wire [511:0] _2825;
    wire [63:0] _2826;
    wire [511:0] _2828;
    wire [383:0] _2829;
    wire [511:0] _2846;
    wire [351:0] _2847;
    wire [511:0] _2858;
    wire [191:0] _2859;
    wire [511:0] _2861;
    wire [31:0] _2862;
    wire [511:0] _2864;
    wire [31:0] _2865;
    wire vdd = 1'b1;
    wire [511:0] _14 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire _2;
    wire [511:0] _13 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire _4;
    wire [383:0] _21;
    wire [31:0] _19 = 32'b00000000000000000000000000000001;
    wire [31:0] _18;
    wire [31:0] _20;
    wire [95:0] _17;
    wire [511:0] _22;
    wire _11 = 1'b1;
    wire _6;
    wire _12;
    wire [511:0] _23;
    wire [511:0] _7;
    reg [511:0] _16;
    wire [31:0] _24;
    wire [31:0] _2866;
    wire [511:0] _2912;
    wire [511:0] _9;
    wire [511:0] _2913;

    /* logic */
    assign _2910 = _2864[31:0];
    assign _2909 = _16[31:0];
    assign _2911 = _2909 + _2910;
    assign _2907 = _2864[63:32];
    assign _2906 = _16[63:32];
    assign _2908 = _2906 + _2907;
    assign _2904 = _2864[95:64];
    assign _2903 = _16[95:64];
    assign _2905 = _2903 + _2904;
    assign _2901 = _2864[127:96];
    assign _2900 = _16[127:96];
    assign _2902 = _2900 + _2901;
    assign _2898 = _2864[159:128];
    assign _2897 = _16[159:128];
    assign _2899 = _2897 + _2898;
    assign _2895 = _2864[191:160];
    assign _2894 = _16[191:160];
    assign _2896 = _2894 + _2895;
    assign _2892 = _2864[223:192];
    assign _2891 = _16[223:192];
    assign _2893 = _2891 + _2892;
    assign _2889 = _2864[255:224];
    assign _2888 = _16[255:224];
    assign _2890 = _2888 + _2889;
    assign _2886 = _2864[287:256];
    assign _2885 = _16[287:256];
    assign _2887 = _2885 + _2886;
    assign _2883 = _2864[319:288];
    assign _2882 = _16[319:288];
    assign _2884 = _2882 + _2883;
    assign _2880 = _2864[351:320];
    assign _2879 = _16[351:320];
    assign _2881 = _2879 + _2880;
    assign _2877 = _2864[383:352];
    assign _2876 = _16[383:352];
    assign _2878 = _2876 + _2877;
    assign _2874 = _2864[415:384];
    assign _2873 = _16[415:384];
    assign _2875 = _2873 + _2874;
    assign _2871 = _2864[447:416];
    assign _2870 = _16[447:416];
    assign _2872 = _2870 + _2871;
    assign _2868 = _2864[479:448];
    assign _2867 = _16[479:448];
    assign _2869 = _2867 + _2868;
    assign _2863 = _2861[447:0];
    assign _2860 = _2858[287:0];
    assign _2857 = _2846[127:0];
    assign _2855 = _2853[31:25];
    assign _2850 = _2848[31:24];
    assign _2848 = _2838 ^ _2844;
    assign _2849 = _2848[23:0];
    assign _2851 = { _2849, _2850 };
    assign _2852 = _2839 + _2851;
    assign _2853 = _2843 ^ _2852;
    assign _2854 = _2853[24:0];
    assign _2856 = { _2854, _2855 };
    assign _2845 = _2828[95:0];
    assign _2842 = _2840[31:20];
    assign _2837 = _2835[31:16];
    assign _2834 = _2828[479:448];
    assign _2835 = _2834 ^ _2832;
    assign _2836 = _2835[15:0];
    assign _2838 = { _2836, _2837 };
    assign _2833 = _2828[319:288];
    assign _2839 = _2833 + _2838;
    assign _2840 = _2831 ^ _2839;
    assign _2841 = _2840[19:0];
    assign _2843 = { _2841, _2842 };
    assign _2831 = _2828[159:128];
    assign _2830 = _2828[127:96];
    assign _2832 = _2830 + _2831;
    assign _2844 = _2832 + _2843;
    assign _2827 = _2825[415:0];
    assign _2824 = _2822[255:0];
    assign _2821 = _2810[223:0];
    assign _2819 = _2817[31:25];
    assign _2814 = _2812[31:24];
    assign _2812 = _2802 ^ _2808;
    assign _2813 = _2812[23:0];
    assign _2815 = { _2813, _2814 };
    assign _2816 = _2803 + _2815;
    assign _2817 = _2807 ^ _2816;
    assign _2818 = _2817[24:0];
    assign _2820 = { _2818, _2819 };
    assign _2809 = _2792[63:0];
    assign _2806 = _2804[31:20];
    assign _2801 = _2799[31:16];
    assign _2798 = _2792[447:416];
    assign _2799 = _2798 ^ _2796;
    assign _2800 = _2799[15:0];
    assign _2802 = { _2800, _2801 };
    assign _2797 = _2792[287:256];
    assign _2803 = _2797 + _2802;
    assign _2804 = _2795 ^ _2803;
    assign _2805 = _2804[19:0];
    assign _2807 = { _2805, _2806 };
    assign _2795 = _2792[255:224];
    assign _2794 = _2792[95:64];
    assign _2796 = _2794 + _2795;
    assign _2808 = _2796 + _2807;
    assign _2791 = _2789[383:0];
    assign _2788 = _2786[351:0];
    assign _2785 = _2774[191:0];
    assign _2783 = _2781[31:25];
    assign _2778 = _2776[31:24];
    assign _2776 = _2766 ^ _2772;
    assign _2777 = _2776[23:0];
    assign _2779 = { _2777, _2778 };
    assign _2780 = _2767 + _2779;
    assign _2781 = _2771 ^ _2780;
    assign _2782 = _2781[24:0];
    assign _2784 = { _2782, _2783 };
    assign _2773 = _2756[31:0];
    assign _2770 = _2768[31:20];
    assign _2765 = _2763[31:16];
    assign _2762 = _2756[415:384];
    assign _2763 = _2762 ^ _2760;
    assign _2764 = _2763[15:0];
    assign _2766 = { _2764, _2765 };
    assign _2761 = _2756[383:352];
    assign _2767 = _2761 + _2766;
    assign _2768 = _2759 ^ _2767;
    assign _2769 = _2768[19:0];
    assign _2771 = { _2769, _2770 };
    assign _2759 = _2756[223:192];
    assign _2758 = _2756[63:32];
    assign _2760 = _2758 + _2759;
    assign _2772 = _2760 + _2771;
    assign _2753 = _2751[319:0];
    assign _2750 = _2743[159:0];
    assign _2748 = _2746[31:25];
    assign _2745 = _2732 + _2741;
    assign _2746 = _2736 ^ _2745;
    assign _2747 = _2746[24:0];
    assign _2749 = { _2747, _2748 };
    assign _2742 = _2722[511:32];
    assign _2743 = { _2742, _2737 };
    assign _2744 = _2743[511:192];
    assign _2751 = { _2744, _2749, _2750 };
    assign _2752 = _2751[511:352];
    assign _2754 = { _2752, _2745, _2753 };
    assign _2755 = _2754[479:0];
    assign _2740 = _2738[31:24];
    assign _2735 = _2733[31:20];
    assign _2731 = _2722[351:320];
    assign _2732 = _2731 + _2730;
    assign _2733 = _2725 ^ _2732;
    assign _2734 = _2733[19:0];
    assign _2736 = { _2734, _2735 };
    assign _2737 = _2726 + _2736;
    assign _2729 = _2727[31:16];
    assign _2725 = _2722[191:160];
    assign _2724 = _2722[31:0];
    assign _2726 = _2724 + _2725;
    assign _2719 = _2717[351:0];
    assign _2716 = _2709[223:0];
    assign _2714 = _2712[31:25];
    assign _2711 = _2697 + _2706;
    assign _2712 = _2701 ^ _2711;
    assign _2713 = _2712[24:0];
    assign _2715 = { _2713, _2714 };
    assign _2708 = _2687[95:0];
    assign _2707 = _2687[511:128];
    assign _2709 = { _2707, _2702, _2708 };
    assign _2710 = _2709[511:256];
    assign _2717 = { _2710, _2715, _2716 };
    assign _2718 = _2717[511:384];
    assign _2720 = { _2718, _2711, _2719 };
    assign _2721 = _2720[479:0];
    assign _2705 = _2703[31:24];
    assign _2700 = _2698[31:20];
    assign _2696 = _2687[383:352];
    assign _2697 = _2696 + _2695;
    assign _2698 = _2690 ^ _2697;
    assign _2699 = _2698[19:0];
    assign _2701 = { _2699, _2700 };
    assign _2702 = _2691 + _2701;
    assign _2694 = _2692[31:16];
    assign _2690 = _2687[255:224];
    assign _2689 = _2687[127:96];
    assign _2691 = _2689 + _2690;
    assign _2686 = _2684[447:0];
    assign _2683 = _2681[319:0];
    assign _2680 = _2669[191:0];
    assign _2678 = _2676[31:25];
    assign _2673 = _2671[31:24];
    assign _2671 = _2661 ^ _2667;
    assign _2672 = _2671[23:0];
    assign _2674 = { _2672, _2673 };
    assign _2675 = _2662 + _2674;
    assign _2676 = _2666 ^ _2675;
    assign _2677 = _2676[24:0];
    assign _2679 = { _2677, _2678 };
    assign _2668 = _2651[63:0];
    assign _2665 = _2663[31:20];
    assign _2660 = _2658[31:16];
    assign _2657 = _2651[479:448];
    assign _2658 = _2657 ^ _2655;
    assign _2659 = _2658[15:0];
    assign _2661 = { _2659, _2660 };
    assign _2656 = _2651[351:320];
    assign _2662 = _2656 + _2661;
    assign _2663 = _2654 ^ _2662;
    assign _2664 = _2663[19:0];
    assign _2666 = { _2664, _2665 };
    assign _2654 = _2651[223:192];
    assign _2653 = _2651[95:64];
    assign _2655 = _2653 + _2654;
    assign _2667 = _2655 + _2666;
    assign _2650 = _2648[415:0];
    assign _2647 = _2645[287:0];
    assign _2644 = _2633[159:0];
    assign _2642 = _2640[31:25];
    assign _2637 = _2635[31:24];
    assign _2635 = _2625 ^ _2631;
    assign _2636 = _2635[23:0];
    assign _2638 = { _2636, _2637 };
    assign _2639 = _2626 + _2638;
    assign _2640 = _2630 ^ _2639;
    assign _2641 = _2640[24:0];
    assign _2643 = { _2641, _2642 };
    assign _2632 = _2615[31:0];
    assign _2629 = _2627[31:20];
    assign _2624 = _2622[31:16];
    assign _2621 = _2615[447:416];
    assign _2622 = _2621 ^ _2619;
    assign _2623 = _2622[15:0];
    assign _2625 = { _2623, _2624 };
    assign _2620 = _2615[319:288];
    assign _2626 = _2620 + _2625;
    assign _2627 = _2618 ^ _2626;
    assign _2628 = _2627[19:0];
    assign _2630 = { _2628, _2629 };
    assign _2618 = _2615[191:160];
    assign _2617 = _2615[63:32];
    assign _2619 = _2617 + _2618;
    assign _2631 = _2619 + _2630;
    assign _2614 = _2612[383:0];
    assign _2611 = _2609[255:0];
    assign _2608 = _2597[127:0];
    assign _2606 = _2604[31:25];
    assign _2601 = _2599[31:24];
    assign _2599 = _2590 ^ _2596;
    assign _2600 = _2599[23:0];
    assign _2602 = { _2600, _2601 };
    assign _2603 = _2591 + _2602;
    assign _2604 = _2595 ^ _2603;
    assign _2605 = _2604[24:0];
    assign _2607 = { _2605, _2606 };
    assign _2594 = _2592[31:20];
    assign _2589 = _2587[31:16];
    assign _2586 = _2580[415:384];
    assign _2587 = _2586 ^ _2584;
    assign _2588 = _2587[15:0];
    assign _2590 = { _2588, _2589 };
    assign _2585 = _2580[287:256];
    assign _2591 = _2585 + _2590;
    assign _2592 = _2583 ^ _2591;
    assign _2593 = _2592[19:0];
    assign _2595 = { _2593, _2594 };
    assign _2583 = _2580[159:128];
    assign _2582 = _2580[31:0];
    assign _2584 = _2582 + _2583;
    assign _2596 = _2584 + _2595;
    assign _2579 = _2577[447:0];
    assign _2576 = _2574[287:0];
    assign _2573 = _2562[127:0];
    assign _2571 = _2569[31:25];
    assign _2566 = _2564[31:24];
    assign _2564 = _2554 ^ _2560;
    assign _2565 = _2564[23:0];
    assign _2567 = { _2565, _2566 };
    assign _2568 = _2555 + _2567;
    assign _2569 = _2559 ^ _2568;
    assign _2570 = _2569[24:0];
    assign _2572 = { _2570, _2571 };
    assign _2561 = _2544[95:0];
    assign _2558 = _2556[31:20];
    assign _2553 = _2551[31:16];
    assign _2550 = _2544[479:448];
    assign _2551 = _2550 ^ _2548;
    assign _2552 = _2551[15:0];
    assign _2554 = { _2552, _2553 };
    assign _2549 = _2544[319:288];
    assign _2555 = _2549 + _2554;
    assign _2556 = _2547 ^ _2555;
    assign _2557 = _2556[19:0];
    assign _2559 = { _2557, _2558 };
    assign _2547 = _2544[159:128];
    assign _2546 = _2544[127:96];
    assign _2548 = _2546 + _2547;
    assign _2560 = _2548 + _2559;
    assign _2543 = _2541[415:0];
    assign _2540 = _2538[255:0];
    assign _2537 = _2526[223:0];
    assign _2535 = _2533[31:25];
    assign _2530 = _2528[31:24];
    assign _2528 = _2518 ^ _2524;
    assign _2529 = _2528[23:0];
    assign _2531 = { _2529, _2530 };
    assign _2532 = _2519 + _2531;
    assign _2533 = _2523 ^ _2532;
    assign _2534 = _2533[24:0];
    assign _2536 = { _2534, _2535 };
    assign _2525 = _2508[63:0];
    assign _2522 = _2520[31:20];
    assign _2517 = _2515[31:16];
    assign _2514 = _2508[447:416];
    assign _2515 = _2514 ^ _2512;
    assign _2516 = _2515[15:0];
    assign _2518 = { _2516, _2517 };
    assign _2513 = _2508[287:256];
    assign _2519 = _2513 + _2518;
    assign _2520 = _2511 ^ _2519;
    assign _2521 = _2520[19:0];
    assign _2523 = { _2521, _2522 };
    assign _2511 = _2508[255:224];
    assign _2510 = _2508[95:64];
    assign _2512 = _2510 + _2511;
    assign _2524 = _2512 + _2523;
    assign _2507 = _2505[383:0];
    assign _2504 = _2502[351:0];
    assign _2501 = _2490[191:0];
    assign _2499 = _2497[31:25];
    assign _2494 = _2492[31:24];
    assign _2492 = _2482 ^ _2488;
    assign _2493 = _2492[23:0];
    assign _2495 = { _2493, _2494 };
    assign _2496 = _2483 + _2495;
    assign _2497 = _2487 ^ _2496;
    assign _2498 = _2497[24:0];
    assign _2500 = { _2498, _2499 };
    assign _2489 = _2472[31:0];
    assign _2486 = _2484[31:20];
    assign _2481 = _2479[31:16];
    assign _2478 = _2472[415:384];
    assign _2479 = _2478 ^ _2476;
    assign _2480 = _2479[15:0];
    assign _2482 = { _2480, _2481 };
    assign _2477 = _2472[383:352];
    assign _2483 = _2477 + _2482;
    assign _2484 = _2475 ^ _2483;
    assign _2485 = _2484[19:0];
    assign _2487 = { _2485, _2486 };
    assign _2475 = _2472[223:192];
    assign _2474 = _2472[63:32];
    assign _2476 = _2474 + _2475;
    assign _2488 = _2476 + _2487;
    assign _2469 = _2467[319:0];
    assign _2466 = _2459[159:0];
    assign _2464 = _2462[31:25];
    assign _2461 = _2448 + _2457;
    assign _2462 = _2452 ^ _2461;
    assign _2463 = _2462[24:0];
    assign _2465 = { _2463, _2464 };
    assign _2458 = _2438[511:32];
    assign _2459 = { _2458, _2453 };
    assign _2460 = _2459[511:192];
    assign _2467 = { _2460, _2465, _2466 };
    assign _2468 = _2467[511:352];
    assign _2470 = { _2468, _2461, _2469 };
    assign _2471 = _2470[479:0];
    assign _2456 = _2454[31:24];
    assign _2451 = _2449[31:20];
    assign _2447 = _2438[351:320];
    assign _2448 = _2447 + _2446;
    assign _2449 = _2441 ^ _2448;
    assign _2450 = _2449[19:0];
    assign _2452 = { _2450, _2451 };
    assign _2453 = _2442 + _2452;
    assign _2445 = _2443[31:16];
    assign _2441 = _2438[191:160];
    assign _2440 = _2438[31:0];
    assign _2442 = _2440 + _2441;
    assign _2435 = _2433[351:0];
    assign _2432 = _2425[223:0];
    assign _2430 = _2428[31:25];
    assign _2427 = _2413 + _2422;
    assign _2428 = _2417 ^ _2427;
    assign _2429 = _2428[24:0];
    assign _2431 = { _2429, _2430 };
    assign _2424 = _2403[95:0];
    assign _2423 = _2403[511:128];
    assign _2425 = { _2423, _2418, _2424 };
    assign _2426 = _2425[511:256];
    assign _2433 = { _2426, _2431, _2432 };
    assign _2434 = _2433[511:384];
    assign _2436 = { _2434, _2427, _2435 };
    assign _2437 = _2436[479:0];
    assign _2421 = _2419[31:24];
    assign _2416 = _2414[31:20];
    assign _2412 = _2403[383:352];
    assign _2413 = _2412 + _2411;
    assign _2414 = _2406 ^ _2413;
    assign _2415 = _2414[19:0];
    assign _2417 = { _2415, _2416 };
    assign _2418 = _2407 + _2417;
    assign _2410 = _2408[31:16];
    assign _2406 = _2403[255:224];
    assign _2405 = _2403[127:96];
    assign _2407 = _2405 + _2406;
    assign _2402 = _2400[447:0];
    assign _2399 = _2397[319:0];
    assign _2396 = _2385[191:0];
    assign _2394 = _2392[31:25];
    assign _2389 = _2387[31:24];
    assign _2387 = _2377 ^ _2383;
    assign _2388 = _2387[23:0];
    assign _2390 = { _2388, _2389 };
    assign _2391 = _2378 + _2390;
    assign _2392 = _2382 ^ _2391;
    assign _2393 = _2392[24:0];
    assign _2395 = { _2393, _2394 };
    assign _2384 = _2367[63:0];
    assign _2381 = _2379[31:20];
    assign _2376 = _2374[31:16];
    assign _2373 = _2367[479:448];
    assign _2374 = _2373 ^ _2371;
    assign _2375 = _2374[15:0];
    assign _2377 = { _2375, _2376 };
    assign _2372 = _2367[351:320];
    assign _2378 = _2372 + _2377;
    assign _2379 = _2370 ^ _2378;
    assign _2380 = _2379[19:0];
    assign _2382 = { _2380, _2381 };
    assign _2370 = _2367[223:192];
    assign _2369 = _2367[95:64];
    assign _2371 = _2369 + _2370;
    assign _2383 = _2371 + _2382;
    assign _2366 = _2364[415:0];
    assign _2363 = _2361[287:0];
    assign _2360 = _2349[159:0];
    assign _2358 = _2356[31:25];
    assign _2353 = _2351[31:24];
    assign _2351 = _2341 ^ _2347;
    assign _2352 = _2351[23:0];
    assign _2354 = { _2352, _2353 };
    assign _2355 = _2342 + _2354;
    assign _2356 = _2346 ^ _2355;
    assign _2357 = _2356[24:0];
    assign _2359 = { _2357, _2358 };
    assign _2348 = _2331[31:0];
    assign _2345 = _2343[31:20];
    assign _2340 = _2338[31:16];
    assign _2337 = _2331[447:416];
    assign _2338 = _2337 ^ _2335;
    assign _2339 = _2338[15:0];
    assign _2341 = { _2339, _2340 };
    assign _2336 = _2331[319:288];
    assign _2342 = _2336 + _2341;
    assign _2343 = _2334 ^ _2342;
    assign _2344 = _2343[19:0];
    assign _2346 = { _2344, _2345 };
    assign _2334 = _2331[191:160];
    assign _2333 = _2331[63:32];
    assign _2335 = _2333 + _2334;
    assign _2347 = _2335 + _2346;
    assign _2330 = _2328[383:0];
    assign _2327 = _2325[255:0];
    assign _2324 = _2313[127:0];
    assign _2322 = _2320[31:25];
    assign _2317 = _2315[31:24];
    assign _2315 = _2306 ^ _2312;
    assign _2316 = _2315[23:0];
    assign _2318 = { _2316, _2317 };
    assign _2319 = _2307 + _2318;
    assign _2320 = _2311 ^ _2319;
    assign _2321 = _2320[24:0];
    assign _2323 = { _2321, _2322 };
    assign _2310 = _2308[31:20];
    assign _2305 = _2303[31:16];
    assign _2302 = _2296[415:384];
    assign _2303 = _2302 ^ _2300;
    assign _2304 = _2303[15:0];
    assign _2306 = { _2304, _2305 };
    assign _2301 = _2296[287:256];
    assign _2307 = _2301 + _2306;
    assign _2308 = _2299 ^ _2307;
    assign _2309 = _2308[19:0];
    assign _2311 = { _2309, _2310 };
    assign _2299 = _2296[159:128];
    assign _2298 = _2296[31:0];
    assign _2300 = _2298 + _2299;
    assign _2312 = _2300 + _2311;
    assign _2295 = _2293[447:0];
    assign _2292 = _2290[287:0];
    assign _2289 = _2278[127:0];
    assign _2287 = _2285[31:25];
    assign _2282 = _2280[31:24];
    assign _2280 = _2270 ^ _2276;
    assign _2281 = _2280[23:0];
    assign _2283 = { _2281, _2282 };
    assign _2284 = _2271 + _2283;
    assign _2285 = _2275 ^ _2284;
    assign _2286 = _2285[24:0];
    assign _2288 = { _2286, _2287 };
    assign _2277 = _2260[95:0];
    assign _2274 = _2272[31:20];
    assign _2269 = _2267[31:16];
    assign _2266 = _2260[479:448];
    assign _2267 = _2266 ^ _2264;
    assign _2268 = _2267[15:0];
    assign _2270 = { _2268, _2269 };
    assign _2265 = _2260[319:288];
    assign _2271 = _2265 + _2270;
    assign _2272 = _2263 ^ _2271;
    assign _2273 = _2272[19:0];
    assign _2275 = { _2273, _2274 };
    assign _2263 = _2260[159:128];
    assign _2262 = _2260[127:96];
    assign _2264 = _2262 + _2263;
    assign _2276 = _2264 + _2275;
    assign _2259 = _2257[415:0];
    assign _2256 = _2254[255:0];
    assign _2253 = _2242[223:0];
    assign _2251 = _2249[31:25];
    assign _2246 = _2244[31:24];
    assign _2244 = _2234 ^ _2240;
    assign _2245 = _2244[23:0];
    assign _2247 = { _2245, _2246 };
    assign _2248 = _2235 + _2247;
    assign _2249 = _2239 ^ _2248;
    assign _2250 = _2249[24:0];
    assign _2252 = { _2250, _2251 };
    assign _2241 = _2224[63:0];
    assign _2238 = _2236[31:20];
    assign _2233 = _2231[31:16];
    assign _2230 = _2224[447:416];
    assign _2231 = _2230 ^ _2228;
    assign _2232 = _2231[15:0];
    assign _2234 = { _2232, _2233 };
    assign _2229 = _2224[287:256];
    assign _2235 = _2229 + _2234;
    assign _2236 = _2227 ^ _2235;
    assign _2237 = _2236[19:0];
    assign _2239 = { _2237, _2238 };
    assign _2227 = _2224[255:224];
    assign _2226 = _2224[95:64];
    assign _2228 = _2226 + _2227;
    assign _2240 = _2228 + _2239;
    assign _2223 = _2221[383:0];
    assign _2220 = _2218[351:0];
    assign _2217 = _2206[191:0];
    assign _2215 = _2213[31:25];
    assign _2210 = _2208[31:24];
    assign _2208 = _2198 ^ _2204;
    assign _2209 = _2208[23:0];
    assign _2211 = { _2209, _2210 };
    assign _2212 = _2199 + _2211;
    assign _2213 = _2203 ^ _2212;
    assign _2214 = _2213[24:0];
    assign _2216 = { _2214, _2215 };
    assign _2205 = _2188[31:0];
    assign _2202 = _2200[31:20];
    assign _2197 = _2195[31:16];
    assign _2194 = _2188[415:384];
    assign _2195 = _2194 ^ _2192;
    assign _2196 = _2195[15:0];
    assign _2198 = { _2196, _2197 };
    assign _2193 = _2188[383:352];
    assign _2199 = _2193 + _2198;
    assign _2200 = _2191 ^ _2199;
    assign _2201 = _2200[19:0];
    assign _2203 = { _2201, _2202 };
    assign _2191 = _2188[223:192];
    assign _2190 = _2188[63:32];
    assign _2192 = _2190 + _2191;
    assign _2204 = _2192 + _2203;
    assign _2185 = _2183[319:0];
    assign _2182 = _2175[159:0];
    assign _2180 = _2178[31:25];
    assign _2177 = _2164 + _2173;
    assign _2178 = _2168 ^ _2177;
    assign _2179 = _2178[24:0];
    assign _2181 = { _2179, _2180 };
    assign _2174 = _2154[511:32];
    assign _2175 = { _2174, _2169 };
    assign _2176 = _2175[511:192];
    assign _2183 = { _2176, _2181, _2182 };
    assign _2184 = _2183[511:352];
    assign _2186 = { _2184, _2177, _2185 };
    assign _2187 = _2186[479:0];
    assign _2172 = _2170[31:24];
    assign _2167 = _2165[31:20];
    assign _2163 = _2154[351:320];
    assign _2164 = _2163 + _2162;
    assign _2165 = _2157 ^ _2164;
    assign _2166 = _2165[19:0];
    assign _2168 = { _2166, _2167 };
    assign _2169 = _2158 + _2168;
    assign _2161 = _2159[31:16];
    assign _2157 = _2154[191:160];
    assign _2156 = _2154[31:0];
    assign _2158 = _2156 + _2157;
    assign _2151 = _2149[351:0];
    assign _2148 = _2141[223:0];
    assign _2146 = _2144[31:25];
    assign _2143 = _2129 + _2138;
    assign _2144 = _2133 ^ _2143;
    assign _2145 = _2144[24:0];
    assign _2147 = { _2145, _2146 };
    assign _2140 = _2119[95:0];
    assign _2139 = _2119[511:128];
    assign _2141 = { _2139, _2134, _2140 };
    assign _2142 = _2141[511:256];
    assign _2149 = { _2142, _2147, _2148 };
    assign _2150 = _2149[511:384];
    assign _2152 = { _2150, _2143, _2151 };
    assign _2153 = _2152[479:0];
    assign _2137 = _2135[31:24];
    assign _2132 = _2130[31:20];
    assign _2128 = _2119[383:352];
    assign _2129 = _2128 + _2127;
    assign _2130 = _2122 ^ _2129;
    assign _2131 = _2130[19:0];
    assign _2133 = { _2131, _2132 };
    assign _2134 = _2123 + _2133;
    assign _2126 = _2124[31:16];
    assign _2122 = _2119[255:224];
    assign _2121 = _2119[127:96];
    assign _2123 = _2121 + _2122;
    assign _2118 = _2116[447:0];
    assign _2115 = _2113[319:0];
    assign _2112 = _2101[191:0];
    assign _2110 = _2108[31:25];
    assign _2105 = _2103[31:24];
    assign _2103 = _2093 ^ _2099;
    assign _2104 = _2103[23:0];
    assign _2106 = { _2104, _2105 };
    assign _2107 = _2094 + _2106;
    assign _2108 = _2098 ^ _2107;
    assign _2109 = _2108[24:0];
    assign _2111 = { _2109, _2110 };
    assign _2100 = _2083[63:0];
    assign _2097 = _2095[31:20];
    assign _2092 = _2090[31:16];
    assign _2089 = _2083[479:448];
    assign _2090 = _2089 ^ _2087;
    assign _2091 = _2090[15:0];
    assign _2093 = { _2091, _2092 };
    assign _2088 = _2083[351:320];
    assign _2094 = _2088 + _2093;
    assign _2095 = _2086 ^ _2094;
    assign _2096 = _2095[19:0];
    assign _2098 = { _2096, _2097 };
    assign _2086 = _2083[223:192];
    assign _2085 = _2083[95:64];
    assign _2087 = _2085 + _2086;
    assign _2099 = _2087 + _2098;
    assign _2082 = _2080[415:0];
    assign _2079 = _2077[287:0];
    assign _2076 = _2065[159:0];
    assign _2074 = _2072[31:25];
    assign _2069 = _2067[31:24];
    assign _2067 = _2057 ^ _2063;
    assign _2068 = _2067[23:0];
    assign _2070 = { _2068, _2069 };
    assign _2071 = _2058 + _2070;
    assign _2072 = _2062 ^ _2071;
    assign _2073 = _2072[24:0];
    assign _2075 = { _2073, _2074 };
    assign _2064 = _2047[31:0];
    assign _2061 = _2059[31:20];
    assign _2056 = _2054[31:16];
    assign _2053 = _2047[447:416];
    assign _2054 = _2053 ^ _2051;
    assign _2055 = _2054[15:0];
    assign _2057 = { _2055, _2056 };
    assign _2052 = _2047[319:288];
    assign _2058 = _2052 + _2057;
    assign _2059 = _2050 ^ _2058;
    assign _2060 = _2059[19:0];
    assign _2062 = { _2060, _2061 };
    assign _2050 = _2047[191:160];
    assign _2049 = _2047[63:32];
    assign _2051 = _2049 + _2050;
    assign _2063 = _2051 + _2062;
    assign _2046 = _2044[383:0];
    assign _2043 = _2041[255:0];
    assign _2040 = _2029[127:0];
    assign _2038 = _2036[31:25];
    assign _2033 = _2031[31:24];
    assign _2031 = _2022 ^ _2028;
    assign _2032 = _2031[23:0];
    assign _2034 = { _2032, _2033 };
    assign _2035 = _2023 + _2034;
    assign _2036 = _2027 ^ _2035;
    assign _2037 = _2036[24:0];
    assign _2039 = { _2037, _2038 };
    assign _2026 = _2024[31:20];
    assign _2021 = _2019[31:16];
    assign _2018 = _2012[415:384];
    assign _2019 = _2018 ^ _2016;
    assign _2020 = _2019[15:0];
    assign _2022 = { _2020, _2021 };
    assign _2017 = _2012[287:256];
    assign _2023 = _2017 + _2022;
    assign _2024 = _2015 ^ _2023;
    assign _2025 = _2024[19:0];
    assign _2027 = { _2025, _2026 };
    assign _2015 = _2012[159:128];
    assign _2014 = _2012[31:0];
    assign _2016 = _2014 + _2015;
    assign _2028 = _2016 + _2027;
    assign _2011 = _2009[447:0];
    assign _2008 = _2006[287:0];
    assign _2005 = _1994[127:0];
    assign _2003 = _2001[31:25];
    assign _1998 = _1996[31:24];
    assign _1996 = _1986 ^ _1992;
    assign _1997 = _1996[23:0];
    assign _1999 = { _1997, _1998 };
    assign _2000 = _1987 + _1999;
    assign _2001 = _1991 ^ _2000;
    assign _2002 = _2001[24:0];
    assign _2004 = { _2002, _2003 };
    assign _1993 = _1976[95:0];
    assign _1990 = _1988[31:20];
    assign _1985 = _1983[31:16];
    assign _1982 = _1976[479:448];
    assign _1983 = _1982 ^ _1980;
    assign _1984 = _1983[15:0];
    assign _1986 = { _1984, _1985 };
    assign _1981 = _1976[319:288];
    assign _1987 = _1981 + _1986;
    assign _1988 = _1979 ^ _1987;
    assign _1989 = _1988[19:0];
    assign _1991 = { _1989, _1990 };
    assign _1979 = _1976[159:128];
    assign _1978 = _1976[127:96];
    assign _1980 = _1978 + _1979;
    assign _1992 = _1980 + _1991;
    assign _1975 = _1973[415:0];
    assign _1972 = _1970[255:0];
    assign _1969 = _1958[223:0];
    assign _1967 = _1965[31:25];
    assign _1962 = _1960[31:24];
    assign _1960 = _1950 ^ _1956;
    assign _1961 = _1960[23:0];
    assign _1963 = { _1961, _1962 };
    assign _1964 = _1951 + _1963;
    assign _1965 = _1955 ^ _1964;
    assign _1966 = _1965[24:0];
    assign _1968 = { _1966, _1967 };
    assign _1957 = _1940[63:0];
    assign _1954 = _1952[31:20];
    assign _1949 = _1947[31:16];
    assign _1946 = _1940[447:416];
    assign _1947 = _1946 ^ _1944;
    assign _1948 = _1947[15:0];
    assign _1950 = { _1948, _1949 };
    assign _1945 = _1940[287:256];
    assign _1951 = _1945 + _1950;
    assign _1952 = _1943 ^ _1951;
    assign _1953 = _1952[19:0];
    assign _1955 = { _1953, _1954 };
    assign _1943 = _1940[255:224];
    assign _1942 = _1940[95:64];
    assign _1944 = _1942 + _1943;
    assign _1956 = _1944 + _1955;
    assign _1939 = _1937[383:0];
    assign _1936 = _1934[351:0];
    assign _1933 = _1922[191:0];
    assign _1931 = _1929[31:25];
    assign _1926 = _1924[31:24];
    assign _1924 = _1914 ^ _1920;
    assign _1925 = _1924[23:0];
    assign _1927 = { _1925, _1926 };
    assign _1928 = _1915 + _1927;
    assign _1929 = _1919 ^ _1928;
    assign _1930 = _1929[24:0];
    assign _1932 = { _1930, _1931 };
    assign _1921 = _1904[31:0];
    assign _1918 = _1916[31:20];
    assign _1913 = _1911[31:16];
    assign _1910 = _1904[415:384];
    assign _1911 = _1910 ^ _1908;
    assign _1912 = _1911[15:0];
    assign _1914 = { _1912, _1913 };
    assign _1909 = _1904[383:352];
    assign _1915 = _1909 + _1914;
    assign _1916 = _1907 ^ _1915;
    assign _1917 = _1916[19:0];
    assign _1919 = { _1917, _1918 };
    assign _1907 = _1904[223:192];
    assign _1906 = _1904[63:32];
    assign _1908 = _1906 + _1907;
    assign _1920 = _1908 + _1919;
    assign _1901 = _1899[319:0];
    assign _1898 = _1891[159:0];
    assign _1896 = _1894[31:25];
    assign _1893 = _1880 + _1889;
    assign _1894 = _1884 ^ _1893;
    assign _1895 = _1894[24:0];
    assign _1897 = { _1895, _1896 };
    assign _1890 = _1870[511:32];
    assign _1891 = { _1890, _1885 };
    assign _1892 = _1891[511:192];
    assign _1899 = { _1892, _1897, _1898 };
    assign _1900 = _1899[511:352];
    assign _1902 = { _1900, _1893, _1901 };
    assign _1903 = _1902[479:0];
    assign _1888 = _1886[31:24];
    assign _1883 = _1881[31:20];
    assign _1879 = _1870[351:320];
    assign _1880 = _1879 + _1878;
    assign _1881 = _1873 ^ _1880;
    assign _1882 = _1881[19:0];
    assign _1884 = { _1882, _1883 };
    assign _1885 = _1874 + _1884;
    assign _1877 = _1875[31:16];
    assign _1873 = _1870[191:160];
    assign _1872 = _1870[31:0];
    assign _1874 = _1872 + _1873;
    assign _1867 = _1865[351:0];
    assign _1864 = _1857[223:0];
    assign _1862 = _1860[31:25];
    assign _1859 = _1845 + _1854;
    assign _1860 = _1849 ^ _1859;
    assign _1861 = _1860[24:0];
    assign _1863 = { _1861, _1862 };
    assign _1856 = _1835[95:0];
    assign _1855 = _1835[511:128];
    assign _1857 = { _1855, _1850, _1856 };
    assign _1858 = _1857[511:256];
    assign _1865 = { _1858, _1863, _1864 };
    assign _1866 = _1865[511:384];
    assign _1868 = { _1866, _1859, _1867 };
    assign _1869 = _1868[479:0];
    assign _1853 = _1851[31:24];
    assign _1848 = _1846[31:20];
    assign _1844 = _1835[383:352];
    assign _1845 = _1844 + _1843;
    assign _1846 = _1838 ^ _1845;
    assign _1847 = _1846[19:0];
    assign _1849 = { _1847, _1848 };
    assign _1850 = _1839 + _1849;
    assign _1842 = _1840[31:16];
    assign _1838 = _1835[255:224];
    assign _1837 = _1835[127:96];
    assign _1839 = _1837 + _1838;
    assign _1834 = _1832[447:0];
    assign _1831 = _1829[319:0];
    assign _1828 = _1817[191:0];
    assign _1826 = _1824[31:25];
    assign _1821 = _1819[31:24];
    assign _1819 = _1809 ^ _1815;
    assign _1820 = _1819[23:0];
    assign _1822 = { _1820, _1821 };
    assign _1823 = _1810 + _1822;
    assign _1824 = _1814 ^ _1823;
    assign _1825 = _1824[24:0];
    assign _1827 = { _1825, _1826 };
    assign _1816 = _1799[63:0];
    assign _1813 = _1811[31:20];
    assign _1808 = _1806[31:16];
    assign _1805 = _1799[479:448];
    assign _1806 = _1805 ^ _1803;
    assign _1807 = _1806[15:0];
    assign _1809 = { _1807, _1808 };
    assign _1804 = _1799[351:320];
    assign _1810 = _1804 + _1809;
    assign _1811 = _1802 ^ _1810;
    assign _1812 = _1811[19:0];
    assign _1814 = { _1812, _1813 };
    assign _1802 = _1799[223:192];
    assign _1801 = _1799[95:64];
    assign _1803 = _1801 + _1802;
    assign _1815 = _1803 + _1814;
    assign _1798 = _1796[415:0];
    assign _1795 = _1793[287:0];
    assign _1792 = _1781[159:0];
    assign _1790 = _1788[31:25];
    assign _1785 = _1783[31:24];
    assign _1783 = _1773 ^ _1779;
    assign _1784 = _1783[23:0];
    assign _1786 = { _1784, _1785 };
    assign _1787 = _1774 + _1786;
    assign _1788 = _1778 ^ _1787;
    assign _1789 = _1788[24:0];
    assign _1791 = { _1789, _1790 };
    assign _1780 = _1763[31:0];
    assign _1777 = _1775[31:20];
    assign _1772 = _1770[31:16];
    assign _1769 = _1763[447:416];
    assign _1770 = _1769 ^ _1767;
    assign _1771 = _1770[15:0];
    assign _1773 = { _1771, _1772 };
    assign _1768 = _1763[319:288];
    assign _1774 = _1768 + _1773;
    assign _1775 = _1766 ^ _1774;
    assign _1776 = _1775[19:0];
    assign _1778 = { _1776, _1777 };
    assign _1766 = _1763[191:160];
    assign _1765 = _1763[63:32];
    assign _1767 = _1765 + _1766;
    assign _1779 = _1767 + _1778;
    assign _1762 = _1760[383:0];
    assign _1759 = _1757[255:0];
    assign _1756 = _1745[127:0];
    assign _1754 = _1752[31:25];
    assign _1749 = _1747[31:24];
    assign _1747 = _1738 ^ _1744;
    assign _1748 = _1747[23:0];
    assign _1750 = { _1748, _1749 };
    assign _1751 = _1739 + _1750;
    assign _1752 = _1743 ^ _1751;
    assign _1753 = _1752[24:0];
    assign _1755 = { _1753, _1754 };
    assign _1742 = _1740[31:20];
    assign _1737 = _1735[31:16];
    assign _1734 = _1728[415:384];
    assign _1735 = _1734 ^ _1732;
    assign _1736 = _1735[15:0];
    assign _1738 = { _1736, _1737 };
    assign _1733 = _1728[287:256];
    assign _1739 = _1733 + _1738;
    assign _1740 = _1731 ^ _1739;
    assign _1741 = _1740[19:0];
    assign _1743 = { _1741, _1742 };
    assign _1731 = _1728[159:128];
    assign _1730 = _1728[31:0];
    assign _1732 = _1730 + _1731;
    assign _1744 = _1732 + _1743;
    assign _1727 = _1725[447:0];
    assign _1724 = _1722[287:0];
    assign _1721 = _1710[127:0];
    assign _1719 = _1717[31:25];
    assign _1714 = _1712[31:24];
    assign _1712 = _1702 ^ _1708;
    assign _1713 = _1712[23:0];
    assign _1715 = { _1713, _1714 };
    assign _1716 = _1703 + _1715;
    assign _1717 = _1707 ^ _1716;
    assign _1718 = _1717[24:0];
    assign _1720 = { _1718, _1719 };
    assign _1709 = _1692[95:0];
    assign _1706 = _1704[31:20];
    assign _1701 = _1699[31:16];
    assign _1698 = _1692[479:448];
    assign _1699 = _1698 ^ _1696;
    assign _1700 = _1699[15:0];
    assign _1702 = { _1700, _1701 };
    assign _1697 = _1692[319:288];
    assign _1703 = _1697 + _1702;
    assign _1704 = _1695 ^ _1703;
    assign _1705 = _1704[19:0];
    assign _1707 = { _1705, _1706 };
    assign _1695 = _1692[159:128];
    assign _1694 = _1692[127:96];
    assign _1696 = _1694 + _1695;
    assign _1708 = _1696 + _1707;
    assign _1691 = _1689[415:0];
    assign _1688 = _1686[255:0];
    assign _1685 = _1674[223:0];
    assign _1683 = _1681[31:25];
    assign _1678 = _1676[31:24];
    assign _1676 = _1666 ^ _1672;
    assign _1677 = _1676[23:0];
    assign _1679 = { _1677, _1678 };
    assign _1680 = _1667 + _1679;
    assign _1681 = _1671 ^ _1680;
    assign _1682 = _1681[24:0];
    assign _1684 = { _1682, _1683 };
    assign _1673 = _1656[63:0];
    assign _1670 = _1668[31:20];
    assign _1665 = _1663[31:16];
    assign _1662 = _1656[447:416];
    assign _1663 = _1662 ^ _1660;
    assign _1664 = _1663[15:0];
    assign _1666 = { _1664, _1665 };
    assign _1661 = _1656[287:256];
    assign _1667 = _1661 + _1666;
    assign _1668 = _1659 ^ _1667;
    assign _1669 = _1668[19:0];
    assign _1671 = { _1669, _1670 };
    assign _1659 = _1656[255:224];
    assign _1658 = _1656[95:64];
    assign _1660 = _1658 + _1659;
    assign _1672 = _1660 + _1671;
    assign _1655 = _1653[383:0];
    assign _1652 = _1650[351:0];
    assign _1649 = _1638[191:0];
    assign _1647 = _1645[31:25];
    assign _1642 = _1640[31:24];
    assign _1640 = _1630 ^ _1636;
    assign _1641 = _1640[23:0];
    assign _1643 = { _1641, _1642 };
    assign _1644 = _1631 + _1643;
    assign _1645 = _1635 ^ _1644;
    assign _1646 = _1645[24:0];
    assign _1648 = { _1646, _1647 };
    assign _1637 = _1620[31:0];
    assign _1634 = _1632[31:20];
    assign _1629 = _1627[31:16];
    assign _1626 = _1620[415:384];
    assign _1627 = _1626 ^ _1624;
    assign _1628 = _1627[15:0];
    assign _1630 = { _1628, _1629 };
    assign _1625 = _1620[383:352];
    assign _1631 = _1625 + _1630;
    assign _1632 = _1623 ^ _1631;
    assign _1633 = _1632[19:0];
    assign _1635 = { _1633, _1634 };
    assign _1623 = _1620[223:192];
    assign _1622 = _1620[63:32];
    assign _1624 = _1622 + _1623;
    assign _1636 = _1624 + _1635;
    assign _1617 = _1615[319:0];
    assign _1614 = _1607[159:0];
    assign _1612 = _1610[31:25];
    assign _1609 = _1596 + _1605;
    assign _1610 = _1600 ^ _1609;
    assign _1611 = _1610[24:0];
    assign _1613 = { _1611, _1612 };
    assign _1606 = _1586[511:32];
    assign _1607 = { _1606, _1601 };
    assign _1608 = _1607[511:192];
    assign _1615 = { _1608, _1613, _1614 };
    assign _1616 = _1615[511:352];
    assign _1618 = { _1616, _1609, _1617 };
    assign _1619 = _1618[479:0];
    assign _1604 = _1602[31:24];
    assign _1599 = _1597[31:20];
    assign _1595 = _1586[351:320];
    assign _1596 = _1595 + _1594;
    assign _1597 = _1589 ^ _1596;
    assign _1598 = _1597[19:0];
    assign _1600 = { _1598, _1599 };
    assign _1601 = _1590 + _1600;
    assign _1593 = _1591[31:16];
    assign _1589 = _1586[191:160];
    assign _1588 = _1586[31:0];
    assign _1590 = _1588 + _1589;
    assign _1583 = _1581[351:0];
    assign _1580 = _1573[223:0];
    assign _1578 = _1576[31:25];
    assign _1575 = _1561 + _1570;
    assign _1576 = _1565 ^ _1575;
    assign _1577 = _1576[24:0];
    assign _1579 = { _1577, _1578 };
    assign _1572 = _1551[95:0];
    assign _1571 = _1551[511:128];
    assign _1573 = { _1571, _1566, _1572 };
    assign _1574 = _1573[511:256];
    assign _1581 = { _1574, _1579, _1580 };
    assign _1582 = _1581[511:384];
    assign _1584 = { _1582, _1575, _1583 };
    assign _1585 = _1584[479:0];
    assign _1569 = _1567[31:24];
    assign _1564 = _1562[31:20];
    assign _1560 = _1551[383:352];
    assign _1561 = _1560 + _1559;
    assign _1562 = _1554 ^ _1561;
    assign _1563 = _1562[19:0];
    assign _1565 = { _1563, _1564 };
    assign _1566 = _1555 + _1565;
    assign _1558 = _1556[31:16];
    assign _1554 = _1551[255:224];
    assign _1553 = _1551[127:96];
    assign _1555 = _1553 + _1554;
    assign _1550 = _1548[447:0];
    assign _1547 = _1545[319:0];
    assign _1544 = _1533[191:0];
    assign _1542 = _1540[31:25];
    assign _1537 = _1535[31:24];
    assign _1535 = _1525 ^ _1531;
    assign _1536 = _1535[23:0];
    assign _1538 = { _1536, _1537 };
    assign _1539 = _1526 + _1538;
    assign _1540 = _1530 ^ _1539;
    assign _1541 = _1540[24:0];
    assign _1543 = { _1541, _1542 };
    assign _1532 = _1515[63:0];
    assign _1529 = _1527[31:20];
    assign _1524 = _1522[31:16];
    assign _1521 = _1515[479:448];
    assign _1522 = _1521 ^ _1519;
    assign _1523 = _1522[15:0];
    assign _1525 = { _1523, _1524 };
    assign _1520 = _1515[351:320];
    assign _1526 = _1520 + _1525;
    assign _1527 = _1518 ^ _1526;
    assign _1528 = _1527[19:0];
    assign _1530 = { _1528, _1529 };
    assign _1518 = _1515[223:192];
    assign _1517 = _1515[95:64];
    assign _1519 = _1517 + _1518;
    assign _1531 = _1519 + _1530;
    assign _1514 = _1512[415:0];
    assign _1511 = _1509[287:0];
    assign _1508 = _1497[159:0];
    assign _1506 = _1504[31:25];
    assign _1501 = _1499[31:24];
    assign _1499 = _1489 ^ _1495;
    assign _1500 = _1499[23:0];
    assign _1502 = { _1500, _1501 };
    assign _1503 = _1490 + _1502;
    assign _1504 = _1494 ^ _1503;
    assign _1505 = _1504[24:0];
    assign _1507 = { _1505, _1506 };
    assign _1496 = _1479[31:0];
    assign _1493 = _1491[31:20];
    assign _1488 = _1486[31:16];
    assign _1485 = _1479[447:416];
    assign _1486 = _1485 ^ _1483;
    assign _1487 = _1486[15:0];
    assign _1489 = { _1487, _1488 };
    assign _1484 = _1479[319:288];
    assign _1490 = _1484 + _1489;
    assign _1491 = _1482 ^ _1490;
    assign _1492 = _1491[19:0];
    assign _1494 = { _1492, _1493 };
    assign _1482 = _1479[191:160];
    assign _1481 = _1479[63:32];
    assign _1483 = _1481 + _1482;
    assign _1495 = _1483 + _1494;
    assign _1478 = _1476[383:0];
    assign _1475 = _1473[255:0];
    assign _1472 = _1461[127:0];
    assign _1470 = _1468[31:25];
    assign _1465 = _1463[31:24];
    assign _1463 = _1454 ^ _1460;
    assign _1464 = _1463[23:0];
    assign _1466 = { _1464, _1465 };
    assign _1467 = _1455 + _1466;
    assign _1468 = _1459 ^ _1467;
    assign _1469 = _1468[24:0];
    assign _1471 = { _1469, _1470 };
    assign _1458 = _1456[31:20];
    assign _1453 = _1451[31:16];
    assign _1450 = _1444[415:384];
    assign _1451 = _1450 ^ _1448;
    assign _1452 = _1451[15:0];
    assign _1454 = { _1452, _1453 };
    assign _1449 = _1444[287:256];
    assign _1455 = _1449 + _1454;
    assign _1456 = _1447 ^ _1455;
    assign _1457 = _1456[19:0];
    assign _1459 = { _1457, _1458 };
    assign _1447 = _1444[159:128];
    assign _1446 = _1444[31:0];
    assign _1448 = _1446 + _1447;
    assign _1460 = _1448 + _1459;
    assign _1443 = _1441[447:0];
    assign _1440 = _1438[287:0];
    assign _1437 = _1426[127:0];
    assign _1435 = _1433[31:25];
    assign _1430 = _1428[31:24];
    assign _1428 = _1418 ^ _1424;
    assign _1429 = _1428[23:0];
    assign _1431 = { _1429, _1430 };
    assign _1432 = _1419 + _1431;
    assign _1433 = _1423 ^ _1432;
    assign _1434 = _1433[24:0];
    assign _1436 = { _1434, _1435 };
    assign _1425 = _1408[95:0];
    assign _1422 = _1420[31:20];
    assign _1417 = _1415[31:16];
    assign _1414 = _1408[479:448];
    assign _1415 = _1414 ^ _1412;
    assign _1416 = _1415[15:0];
    assign _1418 = { _1416, _1417 };
    assign _1413 = _1408[319:288];
    assign _1419 = _1413 + _1418;
    assign _1420 = _1411 ^ _1419;
    assign _1421 = _1420[19:0];
    assign _1423 = { _1421, _1422 };
    assign _1411 = _1408[159:128];
    assign _1410 = _1408[127:96];
    assign _1412 = _1410 + _1411;
    assign _1424 = _1412 + _1423;
    assign _1407 = _1405[415:0];
    assign _1404 = _1402[255:0];
    assign _1401 = _1390[223:0];
    assign _1399 = _1397[31:25];
    assign _1394 = _1392[31:24];
    assign _1392 = _1382 ^ _1388;
    assign _1393 = _1392[23:0];
    assign _1395 = { _1393, _1394 };
    assign _1396 = _1383 + _1395;
    assign _1397 = _1387 ^ _1396;
    assign _1398 = _1397[24:0];
    assign _1400 = { _1398, _1399 };
    assign _1389 = _1372[63:0];
    assign _1386 = _1384[31:20];
    assign _1381 = _1379[31:16];
    assign _1378 = _1372[447:416];
    assign _1379 = _1378 ^ _1376;
    assign _1380 = _1379[15:0];
    assign _1382 = { _1380, _1381 };
    assign _1377 = _1372[287:256];
    assign _1383 = _1377 + _1382;
    assign _1384 = _1375 ^ _1383;
    assign _1385 = _1384[19:0];
    assign _1387 = { _1385, _1386 };
    assign _1375 = _1372[255:224];
    assign _1374 = _1372[95:64];
    assign _1376 = _1374 + _1375;
    assign _1388 = _1376 + _1387;
    assign _1371 = _1369[383:0];
    assign _1368 = _1366[351:0];
    assign _1365 = _1354[191:0];
    assign _1363 = _1361[31:25];
    assign _1358 = _1356[31:24];
    assign _1356 = _1346 ^ _1352;
    assign _1357 = _1356[23:0];
    assign _1359 = { _1357, _1358 };
    assign _1360 = _1347 + _1359;
    assign _1361 = _1351 ^ _1360;
    assign _1362 = _1361[24:0];
    assign _1364 = { _1362, _1363 };
    assign _1353 = _1336[31:0];
    assign _1350 = _1348[31:20];
    assign _1345 = _1343[31:16];
    assign _1342 = _1336[415:384];
    assign _1343 = _1342 ^ _1340;
    assign _1344 = _1343[15:0];
    assign _1346 = { _1344, _1345 };
    assign _1341 = _1336[383:352];
    assign _1347 = _1341 + _1346;
    assign _1348 = _1339 ^ _1347;
    assign _1349 = _1348[19:0];
    assign _1351 = { _1349, _1350 };
    assign _1339 = _1336[223:192];
    assign _1338 = _1336[63:32];
    assign _1340 = _1338 + _1339;
    assign _1352 = _1340 + _1351;
    assign _1333 = _1331[319:0];
    assign _1330 = _1323[159:0];
    assign _1328 = _1326[31:25];
    assign _1325 = _1312 + _1321;
    assign _1326 = _1316 ^ _1325;
    assign _1327 = _1326[24:0];
    assign _1329 = { _1327, _1328 };
    assign _1322 = _1302[511:32];
    assign _1323 = { _1322, _1317 };
    assign _1324 = _1323[511:192];
    assign _1331 = { _1324, _1329, _1330 };
    assign _1332 = _1331[511:352];
    assign _1334 = { _1332, _1325, _1333 };
    assign _1335 = _1334[479:0];
    assign _1320 = _1318[31:24];
    assign _1315 = _1313[31:20];
    assign _1311 = _1302[351:320];
    assign _1312 = _1311 + _1310;
    assign _1313 = _1305 ^ _1312;
    assign _1314 = _1313[19:0];
    assign _1316 = { _1314, _1315 };
    assign _1317 = _1306 + _1316;
    assign _1309 = _1307[31:16];
    assign _1305 = _1302[191:160];
    assign _1304 = _1302[31:0];
    assign _1306 = _1304 + _1305;
    assign _1299 = _1297[351:0];
    assign _1296 = _1289[223:0];
    assign _1294 = _1292[31:25];
    assign _1291 = _1277 + _1286;
    assign _1292 = _1281 ^ _1291;
    assign _1293 = _1292[24:0];
    assign _1295 = { _1293, _1294 };
    assign _1288 = _1267[95:0];
    assign _1287 = _1267[511:128];
    assign _1289 = { _1287, _1282, _1288 };
    assign _1290 = _1289[511:256];
    assign _1297 = { _1290, _1295, _1296 };
    assign _1298 = _1297[511:384];
    assign _1300 = { _1298, _1291, _1299 };
    assign _1301 = _1300[479:0];
    assign _1285 = _1283[31:24];
    assign _1280 = _1278[31:20];
    assign _1276 = _1267[383:352];
    assign _1277 = _1276 + _1275;
    assign _1278 = _1270 ^ _1277;
    assign _1279 = _1278[19:0];
    assign _1281 = { _1279, _1280 };
    assign _1282 = _1271 + _1281;
    assign _1274 = _1272[31:16];
    assign _1270 = _1267[255:224];
    assign _1269 = _1267[127:96];
    assign _1271 = _1269 + _1270;
    assign _1266 = _1264[447:0];
    assign _1263 = _1261[319:0];
    assign _1260 = _1249[191:0];
    assign _1258 = _1256[31:25];
    assign _1253 = _1251[31:24];
    assign _1251 = _1241 ^ _1247;
    assign _1252 = _1251[23:0];
    assign _1254 = { _1252, _1253 };
    assign _1255 = _1242 + _1254;
    assign _1256 = _1246 ^ _1255;
    assign _1257 = _1256[24:0];
    assign _1259 = { _1257, _1258 };
    assign _1248 = _1231[63:0];
    assign _1245 = _1243[31:20];
    assign _1240 = _1238[31:16];
    assign _1237 = _1231[479:448];
    assign _1238 = _1237 ^ _1235;
    assign _1239 = _1238[15:0];
    assign _1241 = { _1239, _1240 };
    assign _1236 = _1231[351:320];
    assign _1242 = _1236 + _1241;
    assign _1243 = _1234 ^ _1242;
    assign _1244 = _1243[19:0];
    assign _1246 = { _1244, _1245 };
    assign _1234 = _1231[223:192];
    assign _1233 = _1231[95:64];
    assign _1235 = _1233 + _1234;
    assign _1247 = _1235 + _1246;
    assign _1230 = _1228[415:0];
    assign _1227 = _1225[287:0];
    assign _1224 = _1213[159:0];
    assign _1222 = _1220[31:25];
    assign _1217 = _1215[31:24];
    assign _1215 = _1205 ^ _1211;
    assign _1216 = _1215[23:0];
    assign _1218 = { _1216, _1217 };
    assign _1219 = _1206 + _1218;
    assign _1220 = _1210 ^ _1219;
    assign _1221 = _1220[24:0];
    assign _1223 = { _1221, _1222 };
    assign _1212 = _1195[31:0];
    assign _1209 = _1207[31:20];
    assign _1204 = _1202[31:16];
    assign _1201 = _1195[447:416];
    assign _1202 = _1201 ^ _1199;
    assign _1203 = _1202[15:0];
    assign _1205 = { _1203, _1204 };
    assign _1200 = _1195[319:288];
    assign _1206 = _1200 + _1205;
    assign _1207 = _1198 ^ _1206;
    assign _1208 = _1207[19:0];
    assign _1210 = { _1208, _1209 };
    assign _1198 = _1195[191:160];
    assign _1197 = _1195[63:32];
    assign _1199 = _1197 + _1198;
    assign _1211 = _1199 + _1210;
    assign _1194 = _1192[383:0];
    assign _1191 = _1189[255:0];
    assign _1188 = _1177[127:0];
    assign _1186 = _1184[31:25];
    assign _1181 = _1179[31:24];
    assign _1179 = _1170 ^ _1176;
    assign _1180 = _1179[23:0];
    assign _1182 = { _1180, _1181 };
    assign _1183 = _1171 + _1182;
    assign _1184 = _1175 ^ _1183;
    assign _1185 = _1184[24:0];
    assign _1187 = { _1185, _1186 };
    assign _1174 = _1172[31:20];
    assign _1169 = _1167[31:16];
    assign _1166 = _1160[415:384];
    assign _1167 = _1166 ^ _1164;
    assign _1168 = _1167[15:0];
    assign _1170 = { _1168, _1169 };
    assign _1165 = _1160[287:256];
    assign _1171 = _1165 + _1170;
    assign _1172 = _1163 ^ _1171;
    assign _1173 = _1172[19:0];
    assign _1175 = { _1173, _1174 };
    assign _1163 = _1160[159:128];
    assign _1162 = _1160[31:0];
    assign _1164 = _1162 + _1163;
    assign _1176 = _1164 + _1175;
    assign _1159 = _1157[447:0];
    assign _1156 = _1154[287:0];
    assign _1153 = _1142[127:0];
    assign _1151 = _1149[31:25];
    assign _1146 = _1144[31:24];
    assign _1144 = _1134 ^ _1140;
    assign _1145 = _1144[23:0];
    assign _1147 = { _1145, _1146 };
    assign _1148 = _1135 + _1147;
    assign _1149 = _1139 ^ _1148;
    assign _1150 = _1149[24:0];
    assign _1152 = { _1150, _1151 };
    assign _1141 = _1124[95:0];
    assign _1138 = _1136[31:20];
    assign _1133 = _1131[31:16];
    assign _1130 = _1124[479:448];
    assign _1131 = _1130 ^ _1128;
    assign _1132 = _1131[15:0];
    assign _1134 = { _1132, _1133 };
    assign _1129 = _1124[319:288];
    assign _1135 = _1129 + _1134;
    assign _1136 = _1127 ^ _1135;
    assign _1137 = _1136[19:0];
    assign _1139 = { _1137, _1138 };
    assign _1127 = _1124[159:128];
    assign _1126 = _1124[127:96];
    assign _1128 = _1126 + _1127;
    assign _1140 = _1128 + _1139;
    assign _1123 = _1121[415:0];
    assign _1120 = _1118[255:0];
    assign _1117 = _1106[223:0];
    assign _1115 = _1113[31:25];
    assign _1110 = _1108[31:24];
    assign _1108 = _1098 ^ _1104;
    assign _1109 = _1108[23:0];
    assign _1111 = { _1109, _1110 };
    assign _1112 = _1099 + _1111;
    assign _1113 = _1103 ^ _1112;
    assign _1114 = _1113[24:0];
    assign _1116 = { _1114, _1115 };
    assign _1105 = _1088[63:0];
    assign _1102 = _1100[31:20];
    assign _1097 = _1095[31:16];
    assign _1094 = _1088[447:416];
    assign _1095 = _1094 ^ _1092;
    assign _1096 = _1095[15:0];
    assign _1098 = { _1096, _1097 };
    assign _1093 = _1088[287:256];
    assign _1099 = _1093 + _1098;
    assign _1100 = _1091 ^ _1099;
    assign _1101 = _1100[19:0];
    assign _1103 = { _1101, _1102 };
    assign _1091 = _1088[255:224];
    assign _1090 = _1088[95:64];
    assign _1092 = _1090 + _1091;
    assign _1104 = _1092 + _1103;
    assign _1087 = _1085[383:0];
    assign _1084 = _1082[351:0];
    assign _1081 = _1070[191:0];
    assign _1079 = _1077[31:25];
    assign _1074 = _1072[31:24];
    assign _1072 = _1062 ^ _1068;
    assign _1073 = _1072[23:0];
    assign _1075 = { _1073, _1074 };
    assign _1076 = _1063 + _1075;
    assign _1077 = _1067 ^ _1076;
    assign _1078 = _1077[24:0];
    assign _1080 = { _1078, _1079 };
    assign _1069 = _1052[31:0];
    assign _1066 = _1064[31:20];
    assign _1061 = _1059[31:16];
    assign _1058 = _1052[415:384];
    assign _1059 = _1058 ^ _1056;
    assign _1060 = _1059[15:0];
    assign _1062 = { _1060, _1061 };
    assign _1057 = _1052[383:352];
    assign _1063 = _1057 + _1062;
    assign _1064 = _1055 ^ _1063;
    assign _1065 = _1064[19:0];
    assign _1067 = { _1065, _1066 };
    assign _1055 = _1052[223:192];
    assign _1054 = _1052[63:32];
    assign _1056 = _1054 + _1055;
    assign _1068 = _1056 + _1067;
    assign _1049 = _1047[319:0];
    assign _1046 = _1039[159:0];
    assign _1044 = _1042[31:25];
    assign _1041 = _1028 + _1037;
    assign _1042 = _1032 ^ _1041;
    assign _1043 = _1042[24:0];
    assign _1045 = { _1043, _1044 };
    assign _1038 = _1018[511:32];
    assign _1039 = { _1038, _1033 };
    assign _1040 = _1039[511:192];
    assign _1047 = { _1040, _1045, _1046 };
    assign _1048 = _1047[511:352];
    assign _1050 = { _1048, _1041, _1049 };
    assign _1051 = _1050[479:0];
    assign _1036 = _1034[31:24];
    assign _1031 = _1029[31:20];
    assign _1027 = _1018[351:320];
    assign _1028 = _1027 + _1026;
    assign _1029 = _1021 ^ _1028;
    assign _1030 = _1029[19:0];
    assign _1032 = { _1030, _1031 };
    assign _1033 = _1022 + _1032;
    assign _1025 = _1023[31:16];
    assign _1021 = _1018[191:160];
    assign _1020 = _1018[31:0];
    assign _1022 = _1020 + _1021;
    assign _1015 = _1013[351:0];
    assign _1012 = _1005[223:0];
    assign _1010 = _1008[31:25];
    assign _1007 = _993 + _1002;
    assign _1008 = _997 ^ _1007;
    assign _1009 = _1008[24:0];
    assign _1011 = { _1009, _1010 };
    assign _1004 = _983[95:0];
    assign _1003 = _983[511:128];
    assign _1005 = { _1003, _998, _1004 };
    assign _1006 = _1005[511:256];
    assign _1013 = { _1006, _1011, _1012 };
    assign _1014 = _1013[511:384];
    assign _1016 = { _1014, _1007, _1015 };
    assign _1017 = _1016[479:0];
    assign _1001 = _999[31:24];
    assign _996 = _994[31:20];
    assign _992 = _983[383:352];
    assign _993 = _992 + _991;
    assign _994 = _986 ^ _993;
    assign _995 = _994[19:0];
    assign _997 = { _995, _996 };
    assign _998 = _987 + _997;
    assign _990 = _988[31:16];
    assign _986 = _983[255:224];
    assign _985 = _983[127:96];
    assign _987 = _985 + _986;
    assign _982 = _980[447:0];
    assign _979 = _977[319:0];
    assign _976 = _965[191:0];
    assign _974 = _972[31:25];
    assign _969 = _967[31:24];
    assign _967 = _957 ^ _963;
    assign _968 = _967[23:0];
    assign _970 = { _968, _969 };
    assign _971 = _958 + _970;
    assign _972 = _962 ^ _971;
    assign _973 = _972[24:0];
    assign _975 = { _973, _974 };
    assign _964 = _947[63:0];
    assign _961 = _959[31:20];
    assign _956 = _954[31:16];
    assign _953 = _947[479:448];
    assign _954 = _953 ^ _951;
    assign _955 = _954[15:0];
    assign _957 = { _955, _956 };
    assign _952 = _947[351:320];
    assign _958 = _952 + _957;
    assign _959 = _950 ^ _958;
    assign _960 = _959[19:0];
    assign _962 = { _960, _961 };
    assign _950 = _947[223:192];
    assign _949 = _947[95:64];
    assign _951 = _949 + _950;
    assign _963 = _951 + _962;
    assign _946 = _944[415:0];
    assign _943 = _941[287:0];
    assign _940 = _929[159:0];
    assign _938 = _936[31:25];
    assign _933 = _931[31:24];
    assign _931 = _921 ^ _927;
    assign _932 = _931[23:0];
    assign _934 = { _932, _933 };
    assign _935 = _922 + _934;
    assign _936 = _926 ^ _935;
    assign _937 = _936[24:0];
    assign _939 = { _937, _938 };
    assign _928 = _911[31:0];
    assign _925 = _923[31:20];
    assign _920 = _918[31:16];
    assign _917 = _911[447:416];
    assign _918 = _917 ^ _915;
    assign _919 = _918[15:0];
    assign _921 = { _919, _920 };
    assign _916 = _911[319:288];
    assign _922 = _916 + _921;
    assign _923 = _914 ^ _922;
    assign _924 = _923[19:0];
    assign _926 = { _924, _925 };
    assign _914 = _911[191:160];
    assign _913 = _911[63:32];
    assign _915 = _913 + _914;
    assign _927 = _915 + _926;
    assign _910 = _908[383:0];
    assign _907 = _905[255:0];
    assign _904 = _893[127:0];
    assign _902 = _900[31:25];
    assign _897 = _895[31:24];
    assign _895 = _886 ^ _892;
    assign _896 = _895[23:0];
    assign _898 = { _896, _897 };
    assign _899 = _887 + _898;
    assign _900 = _891 ^ _899;
    assign _901 = _900[24:0];
    assign _903 = { _901, _902 };
    assign _890 = _888[31:20];
    assign _885 = _883[31:16];
    assign _882 = _876[415:384];
    assign _883 = _882 ^ _880;
    assign _884 = _883[15:0];
    assign _886 = { _884, _885 };
    assign _881 = _876[287:256];
    assign _887 = _881 + _886;
    assign _888 = _879 ^ _887;
    assign _889 = _888[19:0];
    assign _891 = { _889, _890 };
    assign _879 = _876[159:128];
    assign _878 = _876[31:0];
    assign _880 = _878 + _879;
    assign _892 = _880 + _891;
    assign _875 = _873[447:0];
    assign _872 = _870[287:0];
    assign _869 = _858[127:0];
    assign _867 = _865[31:25];
    assign _862 = _860[31:24];
    assign _860 = _850 ^ _856;
    assign _861 = _860[23:0];
    assign _863 = { _861, _862 };
    assign _864 = _851 + _863;
    assign _865 = _855 ^ _864;
    assign _866 = _865[24:0];
    assign _868 = { _866, _867 };
    assign _857 = _840[95:0];
    assign _854 = _852[31:20];
    assign _849 = _847[31:16];
    assign _846 = _840[479:448];
    assign _847 = _846 ^ _844;
    assign _848 = _847[15:0];
    assign _850 = { _848, _849 };
    assign _845 = _840[319:288];
    assign _851 = _845 + _850;
    assign _852 = _843 ^ _851;
    assign _853 = _852[19:0];
    assign _855 = { _853, _854 };
    assign _843 = _840[159:128];
    assign _842 = _840[127:96];
    assign _844 = _842 + _843;
    assign _856 = _844 + _855;
    assign _839 = _837[415:0];
    assign _836 = _834[255:0];
    assign _833 = _822[223:0];
    assign _831 = _829[31:25];
    assign _826 = _824[31:24];
    assign _824 = _814 ^ _820;
    assign _825 = _824[23:0];
    assign _827 = { _825, _826 };
    assign _828 = _815 + _827;
    assign _829 = _819 ^ _828;
    assign _830 = _829[24:0];
    assign _832 = { _830, _831 };
    assign _821 = _804[63:0];
    assign _818 = _816[31:20];
    assign _813 = _811[31:16];
    assign _810 = _804[447:416];
    assign _811 = _810 ^ _808;
    assign _812 = _811[15:0];
    assign _814 = { _812, _813 };
    assign _809 = _804[287:256];
    assign _815 = _809 + _814;
    assign _816 = _807 ^ _815;
    assign _817 = _816[19:0];
    assign _819 = { _817, _818 };
    assign _807 = _804[255:224];
    assign _806 = _804[95:64];
    assign _808 = _806 + _807;
    assign _820 = _808 + _819;
    assign _803 = _801[383:0];
    assign _800 = _798[351:0];
    assign _797 = _786[191:0];
    assign _795 = _793[31:25];
    assign _790 = _788[31:24];
    assign _788 = _778 ^ _784;
    assign _789 = _788[23:0];
    assign _791 = { _789, _790 };
    assign _792 = _779 + _791;
    assign _793 = _783 ^ _792;
    assign _794 = _793[24:0];
    assign _796 = { _794, _795 };
    assign _785 = _768[31:0];
    assign _782 = _780[31:20];
    assign _777 = _775[31:16];
    assign _774 = _768[415:384];
    assign _775 = _774 ^ _772;
    assign _776 = _775[15:0];
    assign _778 = { _776, _777 };
    assign _773 = _768[383:352];
    assign _779 = _773 + _778;
    assign _780 = _771 ^ _779;
    assign _781 = _780[19:0];
    assign _783 = { _781, _782 };
    assign _771 = _768[223:192];
    assign _770 = _768[63:32];
    assign _772 = _770 + _771;
    assign _784 = _772 + _783;
    assign _765 = _763[319:0];
    assign _762 = _755[159:0];
    assign _760 = _758[31:25];
    assign _757 = _744 + _753;
    assign _758 = _748 ^ _757;
    assign _759 = _758[24:0];
    assign _761 = { _759, _760 };
    assign _754 = _734[511:32];
    assign _755 = { _754, _749 };
    assign _756 = _755[511:192];
    assign _763 = { _756, _761, _762 };
    assign _764 = _763[511:352];
    assign _766 = { _764, _757, _765 };
    assign _767 = _766[479:0];
    assign _752 = _750[31:24];
    assign _747 = _745[31:20];
    assign _743 = _734[351:320];
    assign _744 = _743 + _742;
    assign _745 = _737 ^ _744;
    assign _746 = _745[19:0];
    assign _748 = { _746, _747 };
    assign _749 = _738 + _748;
    assign _741 = _739[31:16];
    assign _737 = _734[191:160];
    assign _736 = _734[31:0];
    assign _738 = _736 + _737;
    assign _731 = _729[351:0];
    assign _728 = _721[223:0];
    assign _726 = _724[31:25];
    assign _723 = _709 + _718;
    assign _724 = _713 ^ _723;
    assign _725 = _724[24:0];
    assign _727 = { _725, _726 };
    assign _720 = _699[95:0];
    assign _719 = _699[511:128];
    assign _721 = { _719, _714, _720 };
    assign _722 = _721[511:256];
    assign _729 = { _722, _727, _728 };
    assign _730 = _729[511:384];
    assign _732 = { _730, _723, _731 };
    assign _733 = _732[479:0];
    assign _717 = _715[31:24];
    assign _712 = _710[31:20];
    assign _708 = _699[383:352];
    assign _709 = _708 + _707;
    assign _710 = _702 ^ _709;
    assign _711 = _710[19:0];
    assign _713 = { _711, _712 };
    assign _714 = _703 + _713;
    assign _706 = _704[31:16];
    assign _702 = _699[255:224];
    assign _701 = _699[127:96];
    assign _703 = _701 + _702;
    assign _698 = _696[447:0];
    assign _695 = _693[319:0];
    assign _692 = _681[191:0];
    assign _690 = _688[31:25];
    assign _685 = _683[31:24];
    assign _683 = _673 ^ _679;
    assign _684 = _683[23:0];
    assign _686 = { _684, _685 };
    assign _687 = _674 + _686;
    assign _688 = _678 ^ _687;
    assign _689 = _688[24:0];
    assign _691 = { _689, _690 };
    assign _680 = _663[63:0];
    assign _677 = _675[31:20];
    assign _672 = _670[31:16];
    assign _669 = _663[479:448];
    assign _670 = _669 ^ _667;
    assign _671 = _670[15:0];
    assign _673 = { _671, _672 };
    assign _668 = _663[351:320];
    assign _674 = _668 + _673;
    assign _675 = _666 ^ _674;
    assign _676 = _675[19:0];
    assign _678 = { _676, _677 };
    assign _666 = _663[223:192];
    assign _665 = _663[95:64];
    assign _667 = _665 + _666;
    assign _679 = _667 + _678;
    assign _662 = _660[415:0];
    assign _659 = _657[287:0];
    assign _656 = _645[159:0];
    assign _654 = _652[31:25];
    assign _649 = _647[31:24];
    assign _647 = _637 ^ _643;
    assign _648 = _647[23:0];
    assign _650 = { _648, _649 };
    assign _651 = _638 + _650;
    assign _652 = _642 ^ _651;
    assign _653 = _652[24:0];
    assign _655 = { _653, _654 };
    assign _644 = _627[31:0];
    assign _641 = _639[31:20];
    assign _636 = _634[31:16];
    assign _633 = _627[447:416];
    assign _634 = _633 ^ _631;
    assign _635 = _634[15:0];
    assign _637 = { _635, _636 };
    assign _632 = _627[319:288];
    assign _638 = _632 + _637;
    assign _639 = _630 ^ _638;
    assign _640 = _639[19:0];
    assign _642 = { _640, _641 };
    assign _630 = _627[191:160];
    assign _629 = _627[63:32];
    assign _631 = _629 + _630;
    assign _643 = _631 + _642;
    assign _626 = _624[383:0];
    assign _623 = _621[255:0];
    assign _620 = _609[127:0];
    assign _618 = _616[31:25];
    assign _613 = _611[31:24];
    assign _611 = _602 ^ _608;
    assign _612 = _611[23:0];
    assign _614 = { _612, _613 };
    assign _615 = _603 + _614;
    assign _616 = _607 ^ _615;
    assign _617 = _616[24:0];
    assign _619 = { _617, _618 };
    assign _606 = _604[31:20];
    assign _601 = _599[31:16];
    assign _598 = _592[415:384];
    assign _599 = _598 ^ _596;
    assign _600 = _599[15:0];
    assign _602 = { _600, _601 };
    assign _597 = _592[287:256];
    assign _603 = _597 + _602;
    assign _604 = _595 ^ _603;
    assign _605 = _604[19:0];
    assign _607 = { _605, _606 };
    assign _595 = _592[159:128];
    assign _594 = _592[31:0];
    assign _596 = _594 + _595;
    assign _608 = _596 + _607;
    assign _591 = _589[447:0];
    assign _588 = _586[287:0];
    assign _585 = _574[127:0];
    assign _583 = _581[31:25];
    assign _578 = _576[31:24];
    assign _576 = _566 ^ _572;
    assign _577 = _576[23:0];
    assign _579 = { _577, _578 };
    assign _580 = _567 + _579;
    assign _581 = _571 ^ _580;
    assign _582 = _581[24:0];
    assign _584 = { _582, _583 };
    assign _573 = _556[95:0];
    assign _570 = _568[31:20];
    assign _565 = _563[31:16];
    assign _562 = _556[479:448];
    assign _563 = _562 ^ _560;
    assign _564 = _563[15:0];
    assign _566 = { _564, _565 };
    assign _561 = _556[319:288];
    assign _567 = _561 + _566;
    assign _568 = _559 ^ _567;
    assign _569 = _568[19:0];
    assign _571 = { _569, _570 };
    assign _559 = _556[159:128];
    assign _558 = _556[127:96];
    assign _560 = _558 + _559;
    assign _572 = _560 + _571;
    assign _555 = _553[415:0];
    assign _552 = _550[255:0];
    assign _549 = _538[223:0];
    assign _547 = _545[31:25];
    assign _542 = _540[31:24];
    assign _540 = _530 ^ _536;
    assign _541 = _540[23:0];
    assign _543 = { _541, _542 };
    assign _544 = _531 + _543;
    assign _545 = _535 ^ _544;
    assign _546 = _545[24:0];
    assign _548 = { _546, _547 };
    assign _537 = _520[63:0];
    assign _534 = _532[31:20];
    assign _529 = _527[31:16];
    assign _526 = _520[447:416];
    assign _527 = _526 ^ _524;
    assign _528 = _527[15:0];
    assign _530 = { _528, _529 };
    assign _525 = _520[287:256];
    assign _531 = _525 + _530;
    assign _532 = _523 ^ _531;
    assign _533 = _532[19:0];
    assign _535 = { _533, _534 };
    assign _523 = _520[255:224];
    assign _522 = _520[95:64];
    assign _524 = _522 + _523;
    assign _536 = _524 + _535;
    assign _519 = _517[383:0];
    assign _516 = _514[351:0];
    assign _513 = _502[191:0];
    assign _511 = _509[31:25];
    assign _506 = _504[31:24];
    assign _504 = _494 ^ _500;
    assign _505 = _504[23:0];
    assign _507 = { _505, _506 };
    assign _508 = _495 + _507;
    assign _509 = _499 ^ _508;
    assign _510 = _509[24:0];
    assign _512 = { _510, _511 };
    assign _501 = _484[31:0];
    assign _498 = _496[31:20];
    assign _493 = _491[31:16];
    assign _490 = _484[415:384];
    assign _491 = _490 ^ _488;
    assign _492 = _491[15:0];
    assign _494 = { _492, _493 };
    assign _489 = _484[383:352];
    assign _495 = _489 + _494;
    assign _496 = _487 ^ _495;
    assign _497 = _496[19:0];
    assign _499 = { _497, _498 };
    assign _487 = _484[223:192];
    assign _486 = _484[63:32];
    assign _488 = _486 + _487;
    assign _500 = _488 + _499;
    assign _481 = _479[319:0];
    assign _478 = _471[159:0];
    assign _476 = _474[31:25];
    assign _473 = _460 + _469;
    assign _474 = _464 ^ _473;
    assign _475 = _474[24:0];
    assign _477 = { _475, _476 };
    assign _470 = _450[511:32];
    assign _471 = { _470, _465 };
    assign _472 = _471[511:192];
    assign _479 = { _472, _477, _478 };
    assign _480 = _479[511:352];
    assign _482 = { _480, _473, _481 };
    assign _483 = _482[479:0];
    assign _468 = _466[31:24];
    assign _463 = _461[31:20];
    assign _459 = _450[351:320];
    assign _460 = _459 + _458;
    assign _461 = _453 ^ _460;
    assign _462 = _461[19:0];
    assign _464 = { _462, _463 };
    assign _465 = _454 + _464;
    assign _457 = _455[31:16];
    assign _453 = _450[191:160];
    assign _452 = _450[31:0];
    assign _454 = _452 + _453;
    assign _447 = _445[351:0];
    assign _444 = _437[223:0];
    assign _442 = _440[31:25];
    assign _439 = _425 + _434;
    assign _440 = _429 ^ _439;
    assign _441 = _440[24:0];
    assign _443 = { _441, _442 };
    assign _436 = _415[95:0];
    assign _435 = _415[511:128];
    assign _437 = { _435, _430, _436 };
    assign _438 = _437[511:256];
    assign _445 = { _438, _443, _444 };
    assign _446 = _445[511:384];
    assign _448 = { _446, _439, _447 };
    assign _449 = _448[479:0];
    assign _433 = _431[31:24];
    assign _428 = _426[31:20];
    assign _424 = _415[383:352];
    assign _425 = _424 + _423;
    assign _426 = _418 ^ _425;
    assign _427 = _426[19:0];
    assign _429 = { _427, _428 };
    assign _430 = _419 + _429;
    assign _422 = _420[31:16];
    assign _418 = _415[255:224];
    assign _417 = _415[127:96];
    assign _419 = _417 + _418;
    assign _414 = _412[447:0];
    assign _411 = _409[319:0];
    assign _408 = _397[191:0];
    assign _406 = _404[31:25];
    assign _401 = _399[31:24];
    assign _399 = _389 ^ _395;
    assign _400 = _399[23:0];
    assign _402 = { _400, _401 };
    assign _403 = _390 + _402;
    assign _404 = _394 ^ _403;
    assign _405 = _404[24:0];
    assign _407 = { _405, _406 };
    assign _396 = _379[63:0];
    assign _393 = _391[31:20];
    assign _388 = _386[31:16];
    assign _385 = _379[479:448];
    assign _386 = _385 ^ _383;
    assign _387 = _386[15:0];
    assign _389 = { _387, _388 };
    assign _384 = _379[351:320];
    assign _390 = _384 + _389;
    assign _391 = _382 ^ _390;
    assign _392 = _391[19:0];
    assign _394 = { _392, _393 };
    assign _382 = _379[223:192];
    assign _381 = _379[95:64];
    assign _383 = _381 + _382;
    assign _395 = _383 + _394;
    assign _378 = _376[415:0];
    assign _375 = _373[287:0];
    assign _372 = _361[159:0];
    assign _370 = _368[31:25];
    assign _365 = _363[31:24];
    assign _363 = _353 ^ _359;
    assign _364 = _363[23:0];
    assign _366 = { _364, _365 };
    assign _367 = _354 + _366;
    assign _368 = _358 ^ _367;
    assign _369 = _368[24:0];
    assign _371 = { _369, _370 };
    assign _360 = _343[31:0];
    assign _357 = _355[31:20];
    assign _352 = _350[31:16];
    assign _349 = _343[447:416];
    assign _350 = _349 ^ _347;
    assign _351 = _350[15:0];
    assign _353 = { _351, _352 };
    assign _348 = _343[319:288];
    assign _354 = _348 + _353;
    assign _355 = _346 ^ _354;
    assign _356 = _355[19:0];
    assign _358 = { _356, _357 };
    assign _346 = _343[191:160];
    assign _345 = _343[63:32];
    assign _347 = _345 + _346;
    assign _359 = _347 + _358;
    assign _342 = _340[383:0];
    assign _339 = _337[255:0];
    assign _336 = _325[127:0];
    assign _334 = _332[31:25];
    assign _329 = _327[31:24];
    assign _327 = _318 ^ _324;
    assign _328 = _327[23:0];
    assign _330 = { _328, _329 };
    assign _331 = _319 + _330;
    assign _332 = _323 ^ _331;
    assign _333 = _332[24:0];
    assign _335 = { _333, _334 };
    assign _322 = _320[31:20];
    assign _317 = _315[31:16];
    assign _314 = _308[415:384];
    assign _315 = _314 ^ _312;
    assign _316 = _315[15:0];
    assign _318 = { _316, _317 };
    assign _313 = _308[287:256];
    assign _319 = _313 + _318;
    assign _320 = _311 ^ _319;
    assign _321 = _320[19:0];
    assign _323 = { _321, _322 };
    assign _311 = _308[159:128];
    assign _310 = _308[31:0];
    assign _312 = _310 + _311;
    assign _324 = _312 + _323;
    assign _307 = _305[447:0];
    assign _304 = _302[287:0];
    assign _301 = _290[127:0];
    assign _299 = _297[31:25];
    assign _294 = _292[31:24];
    assign _292 = _282 ^ _288;
    assign _293 = _292[23:0];
    assign _295 = { _293, _294 };
    assign _296 = _283 + _295;
    assign _297 = _287 ^ _296;
    assign _298 = _297[24:0];
    assign _300 = { _298, _299 };
    assign _289 = _272[95:0];
    assign _286 = _284[31:20];
    assign _281 = _279[31:16];
    assign _278 = _272[479:448];
    assign _279 = _278 ^ _276;
    assign _280 = _279[15:0];
    assign _282 = { _280, _281 };
    assign _277 = _272[319:288];
    assign _283 = _277 + _282;
    assign _284 = _275 ^ _283;
    assign _285 = _284[19:0];
    assign _287 = { _285, _286 };
    assign _275 = _272[159:128];
    assign _274 = _272[127:96];
    assign _276 = _274 + _275;
    assign _288 = _276 + _287;
    assign _271 = _269[415:0];
    assign _268 = _266[255:0];
    assign _265 = _254[223:0];
    assign _263 = _261[31:25];
    assign _258 = _256[31:24];
    assign _256 = _246 ^ _252;
    assign _257 = _256[23:0];
    assign _259 = { _257, _258 };
    assign _260 = _247 + _259;
    assign _261 = _251 ^ _260;
    assign _262 = _261[24:0];
    assign _264 = { _262, _263 };
    assign _253 = _236[63:0];
    assign _250 = _248[31:20];
    assign _245 = _243[31:16];
    assign _242 = _236[447:416];
    assign _243 = _242 ^ _240;
    assign _244 = _243[15:0];
    assign _246 = { _244, _245 };
    assign _241 = _236[287:256];
    assign _247 = _241 + _246;
    assign _248 = _239 ^ _247;
    assign _249 = _248[19:0];
    assign _251 = { _249, _250 };
    assign _239 = _236[255:224];
    assign _238 = _236[95:64];
    assign _240 = _238 + _239;
    assign _252 = _240 + _251;
    assign _235 = _233[383:0];
    assign _232 = _230[351:0];
    assign _229 = _218[191:0];
    assign _227 = _225[31:25];
    assign _222 = _220[31:24];
    assign _220 = _210 ^ _216;
    assign _221 = _220[23:0];
    assign _223 = { _221, _222 };
    assign _224 = _211 + _223;
    assign _225 = _215 ^ _224;
    assign _226 = _225[24:0];
    assign _228 = { _226, _227 };
    assign _217 = _200[31:0];
    assign _214 = _212[31:20];
    assign _209 = _207[31:16];
    assign _206 = _200[415:384];
    assign _207 = _206 ^ _204;
    assign _208 = _207[15:0];
    assign _210 = { _208, _209 };
    assign _205 = _200[383:352];
    assign _211 = _205 + _210;
    assign _212 = _203 ^ _211;
    assign _213 = _212[19:0];
    assign _215 = { _213, _214 };
    assign _203 = _200[223:192];
    assign _202 = _200[63:32];
    assign _204 = _202 + _203;
    assign _216 = _204 + _215;
    assign _197 = _195[319:0];
    assign _194 = _187[159:0];
    assign _192 = _190[31:25];
    assign _189 = _176 + _185;
    assign _190 = _180 ^ _189;
    assign _191 = _190[24:0];
    assign _193 = { _191, _192 };
    assign _186 = _166[511:32];
    assign _187 = { _186, _181 };
    assign _188 = _187[511:192];
    assign _195 = { _188, _193, _194 };
    assign _196 = _195[511:352];
    assign _198 = { _196, _189, _197 };
    assign _199 = _198[479:0];
    assign _184 = _182[31:24];
    assign _179 = _177[31:20];
    assign _175 = _166[351:320];
    assign _176 = _175 + _174;
    assign _177 = _169 ^ _176;
    assign _178 = _177[19:0];
    assign _180 = { _178, _179 };
    assign _181 = _170 + _180;
    assign _173 = _171[31:16];
    assign _169 = _166[191:160];
    assign _168 = _166[31:0];
    assign _170 = _168 + _169;
    assign _163 = _161[351:0];
    assign _160 = _153[223:0];
    assign _158 = _156[31:25];
    assign _155 = _141 + _150;
    assign _156 = _145 ^ _155;
    assign _157 = _156[24:0];
    assign _159 = { _157, _158 };
    assign _152 = _131[95:0];
    assign _151 = _131[511:128];
    assign _153 = { _151, _146, _152 };
    assign _154 = _153[511:256];
    assign _161 = { _154, _159, _160 };
    assign _162 = _161[511:384];
    assign _164 = { _162, _155, _163 };
    assign _165 = _164[479:0];
    assign _149 = _147[31:24];
    assign _144 = _142[31:20];
    assign _140 = _131[383:352];
    assign _141 = _140 + _139;
    assign _142 = _134 ^ _141;
    assign _143 = _142[19:0];
    assign _145 = { _143, _144 };
    assign _146 = _135 + _145;
    assign _138 = _136[31:16];
    assign _134 = _131[255:224];
    assign _133 = _131[127:96];
    assign _135 = _133 + _134;
    assign _130 = _128[447:0];
    assign _127 = _125[319:0];
    assign _124 = _113[191:0];
    assign _122 = _120[31:25];
    assign _117 = _115[31:24];
    assign _115 = _105 ^ _111;
    assign _116 = _115[23:0];
    assign _118 = { _116, _117 };
    assign _119 = _106 + _118;
    assign _120 = _110 ^ _119;
    assign _121 = _120[24:0];
    assign _123 = { _121, _122 };
    assign _112 = _95[63:0];
    assign _109 = _107[31:20];
    assign _104 = _102[31:16];
    assign _101 = _95[479:448];
    assign _102 = _101 ^ _99;
    assign _103 = _102[15:0];
    assign _105 = { _103, _104 };
    assign _100 = _95[351:320];
    assign _106 = _100 + _105;
    assign _107 = _98 ^ _106;
    assign _108 = _107[19:0];
    assign _110 = { _108, _109 };
    assign _98 = _95[223:192];
    assign _97 = _95[95:64];
    assign _99 = _97 + _98;
    assign _111 = _99 + _110;
    assign _94 = _92[415:0];
    assign _91 = _89[287:0];
    assign _88 = _77[159:0];
    assign _86 = _84[31:25];
    assign _81 = _79[31:24];
    assign _79 = _69 ^ _75;
    assign _80 = _79[23:0];
    assign _82 = { _80, _81 };
    assign _83 = _70 + _82;
    assign _84 = _74 ^ _83;
    assign _85 = _84[24:0];
    assign _87 = { _85, _86 };
    assign _76 = _59[31:0];
    assign _73 = _71[31:20];
    assign _68 = _66[31:16];
    assign _65 = _59[447:416];
    assign _66 = _65 ^ _63;
    assign _67 = _66[15:0];
    assign _69 = { _67, _68 };
    assign _64 = _59[319:288];
    assign _70 = _64 + _69;
    assign _71 = _62 ^ _70;
    assign _72 = _71[19:0];
    assign _74 = { _72, _73 };
    assign _62 = _59[191:160];
    assign _61 = _59[63:32];
    assign _63 = _61 + _62;
    assign _75 = _63 + _74;
    assign _58 = _56[383:0];
    assign _55 = _53[255:0];
    assign _52 = _41[127:0];
    assign _50 = _48[31:25];
    assign _45 = _43[31:24];
    assign _43 = _34 ^ _40;
    assign _44 = _43[23:0];
    assign _46 = { _44, _45 };
    assign _47 = _35 + _46;
    assign _48 = _39 ^ _47;
    assign _49 = _48[24:0];
    assign _51 = { _49, _50 };
    assign _38 = _36[31:20];
    assign _33 = _31[31:16];
    assign _30 = _16[415:384];
    assign _31 = _30 ^ _28;
    assign _32 = _31[15:0];
    assign _34 = { _32, _33 };
    assign _29 = _16[287:256];
    assign _35 = _29 + _34;
    assign _36 = _27 ^ _35;
    assign _37 = _36[19:0];
    assign _39 = { _37, _38 };
    assign _27 = _16[159:128];
    assign _26 = _16[31:0];
    assign _28 = _26 + _27;
    assign _40 = _28 + _39;
    assign _25 = _16[511:32];
    assign _41 = { _25, _40 };
    assign _42 = _41[511:160];
    assign _53 = { _42, _51, _52 };
    assign _54 = _53[511:288];
    assign _56 = { _54, _47, _55 };
    assign _57 = _56[511:416];
    assign _59 = { _57, _46, _58 };
    assign _60 = _59[511:64];
    assign _77 = { _60, _75, _76 };
    assign _78 = _77[511:192];
    assign _89 = { _78, _87, _88 };
    assign _90 = _89[511:320];
    assign _92 = { _90, _83, _91 };
    assign _93 = _92[511:448];
    assign _95 = { _93, _82, _94 };
    assign _96 = _95[511:96];
    assign _113 = { _96, _111, _112 };
    assign _114 = _113[511:224];
    assign _125 = { _114, _123, _124 };
    assign _126 = _125[511:352];
    assign _128 = { _126, _119, _127 };
    assign _129 = _128[511:480];
    assign _131 = { _129, _118, _130 };
    assign _132 = _131[511:480];
    assign _136 = _132 ^ _135;
    assign _137 = _136[15:0];
    assign _139 = { _137, _138 };
    assign _147 = _139 ^ _146;
    assign _148 = _147[23:0];
    assign _150 = { _148, _149 };
    assign _166 = { _150, _165 };
    assign _167 = _166[511:480];
    assign _171 = _167 ^ _170;
    assign _172 = _171[15:0];
    assign _174 = { _172, _173 };
    assign _182 = _174 ^ _181;
    assign _183 = _182[23:0];
    assign _185 = { _183, _184 };
    assign _200 = { _185, _199 };
    assign _201 = _200[511:64];
    assign _218 = { _201, _216, _217 };
    assign _219 = _218[511:224];
    assign _230 = { _219, _228, _229 };
    assign _231 = _230[511:384];
    assign _233 = { _231, _224, _232 };
    assign _234 = _233[511:416];
    assign _236 = { _234, _223, _235 };
    assign _237 = _236[511:96];
    assign _254 = { _237, _252, _253 };
    assign _255 = _254[511:256];
    assign _266 = { _255, _264, _265 };
    assign _267 = _266[511:288];
    assign _269 = { _267, _260, _268 };
    assign _270 = _269[511:448];
    assign _272 = { _270, _259, _271 };
    assign _273 = _272[511:128];
    assign _290 = { _273, _288, _289 };
    assign _291 = _290[511:160];
    assign _302 = { _291, _300, _301 };
    assign _303 = _302[511:320];
    assign _305 = { _303, _296, _304 };
    assign _306 = _305[511:480];
    assign _308 = { _306, _295, _307 };
    assign _309 = _308[511:32];
    assign _325 = { _309, _324 };
    assign _326 = _325[511:160];
    assign _337 = { _326, _335, _336 };
    assign _338 = _337[511:288];
    assign _340 = { _338, _331, _339 };
    assign _341 = _340[511:416];
    assign _343 = { _341, _330, _342 };
    assign _344 = _343[511:64];
    assign _361 = { _344, _359, _360 };
    assign _362 = _361[511:192];
    assign _373 = { _362, _371, _372 };
    assign _374 = _373[511:320];
    assign _376 = { _374, _367, _375 };
    assign _377 = _376[511:448];
    assign _379 = { _377, _366, _378 };
    assign _380 = _379[511:96];
    assign _397 = { _380, _395, _396 };
    assign _398 = _397[511:224];
    assign _409 = { _398, _407, _408 };
    assign _410 = _409[511:352];
    assign _412 = { _410, _403, _411 };
    assign _413 = _412[511:480];
    assign _415 = { _413, _402, _414 };
    assign _416 = _415[511:480];
    assign _420 = _416 ^ _419;
    assign _421 = _420[15:0];
    assign _423 = { _421, _422 };
    assign _431 = _423 ^ _430;
    assign _432 = _431[23:0];
    assign _434 = { _432, _433 };
    assign _450 = { _434, _449 };
    assign _451 = _450[511:480];
    assign _455 = _451 ^ _454;
    assign _456 = _455[15:0];
    assign _458 = { _456, _457 };
    assign _466 = _458 ^ _465;
    assign _467 = _466[23:0];
    assign _469 = { _467, _468 };
    assign _484 = { _469, _483 };
    assign _485 = _484[511:64];
    assign _502 = { _485, _500, _501 };
    assign _503 = _502[511:224];
    assign _514 = { _503, _512, _513 };
    assign _515 = _514[511:384];
    assign _517 = { _515, _508, _516 };
    assign _518 = _517[511:416];
    assign _520 = { _518, _507, _519 };
    assign _521 = _520[511:96];
    assign _538 = { _521, _536, _537 };
    assign _539 = _538[511:256];
    assign _550 = { _539, _548, _549 };
    assign _551 = _550[511:288];
    assign _553 = { _551, _544, _552 };
    assign _554 = _553[511:448];
    assign _556 = { _554, _543, _555 };
    assign _557 = _556[511:128];
    assign _574 = { _557, _572, _573 };
    assign _575 = _574[511:160];
    assign _586 = { _575, _584, _585 };
    assign _587 = _586[511:320];
    assign _589 = { _587, _580, _588 };
    assign _590 = _589[511:480];
    assign _592 = { _590, _579, _591 };
    assign _593 = _592[511:32];
    assign _609 = { _593, _608 };
    assign _610 = _609[511:160];
    assign _621 = { _610, _619, _620 };
    assign _622 = _621[511:288];
    assign _624 = { _622, _615, _623 };
    assign _625 = _624[511:416];
    assign _627 = { _625, _614, _626 };
    assign _628 = _627[511:64];
    assign _645 = { _628, _643, _644 };
    assign _646 = _645[511:192];
    assign _657 = { _646, _655, _656 };
    assign _658 = _657[511:320];
    assign _660 = { _658, _651, _659 };
    assign _661 = _660[511:448];
    assign _663 = { _661, _650, _662 };
    assign _664 = _663[511:96];
    assign _681 = { _664, _679, _680 };
    assign _682 = _681[511:224];
    assign _693 = { _682, _691, _692 };
    assign _694 = _693[511:352];
    assign _696 = { _694, _687, _695 };
    assign _697 = _696[511:480];
    assign _699 = { _697, _686, _698 };
    assign _700 = _699[511:480];
    assign _704 = _700 ^ _703;
    assign _705 = _704[15:0];
    assign _707 = { _705, _706 };
    assign _715 = _707 ^ _714;
    assign _716 = _715[23:0];
    assign _718 = { _716, _717 };
    assign _734 = { _718, _733 };
    assign _735 = _734[511:480];
    assign _739 = _735 ^ _738;
    assign _740 = _739[15:0];
    assign _742 = { _740, _741 };
    assign _750 = _742 ^ _749;
    assign _751 = _750[23:0];
    assign _753 = { _751, _752 };
    assign _768 = { _753, _767 };
    assign _769 = _768[511:64];
    assign _786 = { _769, _784, _785 };
    assign _787 = _786[511:224];
    assign _798 = { _787, _796, _797 };
    assign _799 = _798[511:384];
    assign _801 = { _799, _792, _800 };
    assign _802 = _801[511:416];
    assign _804 = { _802, _791, _803 };
    assign _805 = _804[511:96];
    assign _822 = { _805, _820, _821 };
    assign _823 = _822[511:256];
    assign _834 = { _823, _832, _833 };
    assign _835 = _834[511:288];
    assign _837 = { _835, _828, _836 };
    assign _838 = _837[511:448];
    assign _840 = { _838, _827, _839 };
    assign _841 = _840[511:128];
    assign _858 = { _841, _856, _857 };
    assign _859 = _858[511:160];
    assign _870 = { _859, _868, _869 };
    assign _871 = _870[511:320];
    assign _873 = { _871, _864, _872 };
    assign _874 = _873[511:480];
    assign _876 = { _874, _863, _875 };
    assign _877 = _876[511:32];
    assign _893 = { _877, _892 };
    assign _894 = _893[511:160];
    assign _905 = { _894, _903, _904 };
    assign _906 = _905[511:288];
    assign _908 = { _906, _899, _907 };
    assign _909 = _908[511:416];
    assign _911 = { _909, _898, _910 };
    assign _912 = _911[511:64];
    assign _929 = { _912, _927, _928 };
    assign _930 = _929[511:192];
    assign _941 = { _930, _939, _940 };
    assign _942 = _941[511:320];
    assign _944 = { _942, _935, _943 };
    assign _945 = _944[511:448];
    assign _947 = { _945, _934, _946 };
    assign _948 = _947[511:96];
    assign _965 = { _948, _963, _964 };
    assign _966 = _965[511:224];
    assign _977 = { _966, _975, _976 };
    assign _978 = _977[511:352];
    assign _980 = { _978, _971, _979 };
    assign _981 = _980[511:480];
    assign _983 = { _981, _970, _982 };
    assign _984 = _983[511:480];
    assign _988 = _984 ^ _987;
    assign _989 = _988[15:0];
    assign _991 = { _989, _990 };
    assign _999 = _991 ^ _998;
    assign _1000 = _999[23:0];
    assign _1002 = { _1000, _1001 };
    assign _1018 = { _1002, _1017 };
    assign _1019 = _1018[511:480];
    assign _1023 = _1019 ^ _1022;
    assign _1024 = _1023[15:0];
    assign _1026 = { _1024, _1025 };
    assign _1034 = _1026 ^ _1033;
    assign _1035 = _1034[23:0];
    assign _1037 = { _1035, _1036 };
    assign _1052 = { _1037, _1051 };
    assign _1053 = _1052[511:64];
    assign _1070 = { _1053, _1068, _1069 };
    assign _1071 = _1070[511:224];
    assign _1082 = { _1071, _1080, _1081 };
    assign _1083 = _1082[511:384];
    assign _1085 = { _1083, _1076, _1084 };
    assign _1086 = _1085[511:416];
    assign _1088 = { _1086, _1075, _1087 };
    assign _1089 = _1088[511:96];
    assign _1106 = { _1089, _1104, _1105 };
    assign _1107 = _1106[511:256];
    assign _1118 = { _1107, _1116, _1117 };
    assign _1119 = _1118[511:288];
    assign _1121 = { _1119, _1112, _1120 };
    assign _1122 = _1121[511:448];
    assign _1124 = { _1122, _1111, _1123 };
    assign _1125 = _1124[511:128];
    assign _1142 = { _1125, _1140, _1141 };
    assign _1143 = _1142[511:160];
    assign _1154 = { _1143, _1152, _1153 };
    assign _1155 = _1154[511:320];
    assign _1157 = { _1155, _1148, _1156 };
    assign _1158 = _1157[511:480];
    assign _1160 = { _1158, _1147, _1159 };
    assign _1161 = _1160[511:32];
    assign _1177 = { _1161, _1176 };
    assign _1178 = _1177[511:160];
    assign _1189 = { _1178, _1187, _1188 };
    assign _1190 = _1189[511:288];
    assign _1192 = { _1190, _1183, _1191 };
    assign _1193 = _1192[511:416];
    assign _1195 = { _1193, _1182, _1194 };
    assign _1196 = _1195[511:64];
    assign _1213 = { _1196, _1211, _1212 };
    assign _1214 = _1213[511:192];
    assign _1225 = { _1214, _1223, _1224 };
    assign _1226 = _1225[511:320];
    assign _1228 = { _1226, _1219, _1227 };
    assign _1229 = _1228[511:448];
    assign _1231 = { _1229, _1218, _1230 };
    assign _1232 = _1231[511:96];
    assign _1249 = { _1232, _1247, _1248 };
    assign _1250 = _1249[511:224];
    assign _1261 = { _1250, _1259, _1260 };
    assign _1262 = _1261[511:352];
    assign _1264 = { _1262, _1255, _1263 };
    assign _1265 = _1264[511:480];
    assign _1267 = { _1265, _1254, _1266 };
    assign _1268 = _1267[511:480];
    assign _1272 = _1268 ^ _1271;
    assign _1273 = _1272[15:0];
    assign _1275 = { _1273, _1274 };
    assign _1283 = _1275 ^ _1282;
    assign _1284 = _1283[23:0];
    assign _1286 = { _1284, _1285 };
    assign _1302 = { _1286, _1301 };
    assign _1303 = _1302[511:480];
    assign _1307 = _1303 ^ _1306;
    assign _1308 = _1307[15:0];
    assign _1310 = { _1308, _1309 };
    assign _1318 = _1310 ^ _1317;
    assign _1319 = _1318[23:0];
    assign _1321 = { _1319, _1320 };
    assign _1336 = { _1321, _1335 };
    assign _1337 = _1336[511:64];
    assign _1354 = { _1337, _1352, _1353 };
    assign _1355 = _1354[511:224];
    assign _1366 = { _1355, _1364, _1365 };
    assign _1367 = _1366[511:384];
    assign _1369 = { _1367, _1360, _1368 };
    assign _1370 = _1369[511:416];
    assign _1372 = { _1370, _1359, _1371 };
    assign _1373 = _1372[511:96];
    assign _1390 = { _1373, _1388, _1389 };
    assign _1391 = _1390[511:256];
    assign _1402 = { _1391, _1400, _1401 };
    assign _1403 = _1402[511:288];
    assign _1405 = { _1403, _1396, _1404 };
    assign _1406 = _1405[511:448];
    assign _1408 = { _1406, _1395, _1407 };
    assign _1409 = _1408[511:128];
    assign _1426 = { _1409, _1424, _1425 };
    assign _1427 = _1426[511:160];
    assign _1438 = { _1427, _1436, _1437 };
    assign _1439 = _1438[511:320];
    assign _1441 = { _1439, _1432, _1440 };
    assign _1442 = _1441[511:480];
    assign _1444 = { _1442, _1431, _1443 };
    assign _1445 = _1444[511:32];
    assign _1461 = { _1445, _1460 };
    assign _1462 = _1461[511:160];
    assign _1473 = { _1462, _1471, _1472 };
    assign _1474 = _1473[511:288];
    assign _1476 = { _1474, _1467, _1475 };
    assign _1477 = _1476[511:416];
    assign _1479 = { _1477, _1466, _1478 };
    assign _1480 = _1479[511:64];
    assign _1497 = { _1480, _1495, _1496 };
    assign _1498 = _1497[511:192];
    assign _1509 = { _1498, _1507, _1508 };
    assign _1510 = _1509[511:320];
    assign _1512 = { _1510, _1503, _1511 };
    assign _1513 = _1512[511:448];
    assign _1515 = { _1513, _1502, _1514 };
    assign _1516 = _1515[511:96];
    assign _1533 = { _1516, _1531, _1532 };
    assign _1534 = _1533[511:224];
    assign _1545 = { _1534, _1543, _1544 };
    assign _1546 = _1545[511:352];
    assign _1548 = { _1546, _1539, _1547 };
    assign _1549 = _1548[511:480];
    assign _1551 = { _1549, _1538, _1550 };
    assign _1552 = _1551[511:480];
    assign _1556 = _1552 ^ _1555;
    assign _1557 = _1556[15:0];
    assign _1559 = { _1557, _1558 };
    assign _1567 = _1559 ^ _1566;
    assign _1568 = _1567[23:0];
    assign _1570 = { _1568, _1569 };
    assign _1586 = { _1570, _1585 };
    assign _1587 = _1586[511:480];
    assign _1591 = _1587 ^ _1590;
    assign _1592 = _1591[15:0];
    assign _1594 = { _1592, _1593 };
    assign _1602 = _1594 ^ _1601;
    assign _1603 = _1602[23:0];
    assign _1605 = { _1603, _1604 };
    assign _1620 = { _1605, _1619 };
    assign _1621 = _1620[511:64];
    assign _1638 = { _1621, _1636, _1637 };
    assign _1639 = _1638[511:224];
    assign _1650 = { _1639, _1648, _1649 };
    assign _1651 = _1650[511:384];
    assign _1653 = { _1651, _1644, _1652 };
    assign _1654 = _1653[511:416];
    assign _1656 = { _1654, _1643, _1655 };
    assign _1657 = _1656[511:96];
    assign _1674 = { _1657, _1672, _1673 };
    assign _1675 = _1674[511:256];
    assign _1686 = { _1675, _1684, _1685 };
    assign _1687 = _1686[511:288];
    assign _1689 = { _1687, _1680, _1688 };
    assign _1690 = _1689[511:448];
    assign _1692 = { _1690, _1679, _1691 };
    assign _1693 = _1692[511:128];
    assign _1710 = { _1693, _1708, _1709 };
    assign _1711 = _1710[511:160];
    assign _1722 = { _1711, _1720, _1721 };
    assign _1723 = _1722[511:320];
    assign _1725 = { _1723, _1716, _1724 };
    assign _1726 = _1725[511:480];
    assign _1728 = { _1726, _1715, _1727 };
    assign _1729 = _1728[511:32];
    assign _1745 = { _1729, _1744 };
    assign _1746 = _1745[511:160];
    assign _1757 = { _1746, _1755, _1756 };
    assign _1758 = _1757[511:288];
    assign _1760 = { _1758, _1751, _1759 };
    assign _1761 = _1760[511:416];
    assign _1763 = { _1761, _1750, _1762 };
    assign _1764 = _1763[511:64];
    assign _1781 = { _1764, _1779, _1780 };
    assign _1782 = _1781[511:192];
    assign _1793 = { _1782, _1791, _1792 };
    assign _1794 = _1793[511:320];
    assign _1796 = { _1794, _1787, _1795 };
    assign _1797 = _1796[511:448];
    assign _1799 = { _1797, _1786, _1798 };
    assign _1800 = _1799[511:96];
    assign _1817 = { _1800, _1815, _1816 };
    assign _1818 = _1817[511:224];
    assign _1829 = { _1818, _1827, _1828 };
    assign _1830 = _1829[511:352];
    assign _1832 = { _1830, _1823, _1831 };
    assign _1833 = _1832[511:480];
    assign _1835 = { _1833, _1822, _1834 };
    assign _1836 = _1835[511:480];
    assign _1840 = _1836 ^ _1839;
    assign _1841 = _1840[15:0];
    assign _1843 = { _1841, _1842 };
    assign _1851 = _1843 ^ _1850;
    assign _1852 = _1851[23:0];
    assign _1854 = { _1852, _1853 };
    assign _1870 = { _1854, _1869 };
    assign _1871 = _1870[511:480];
    assign _1875 = _1871 ^ _1874;
    assign _1876 = _1875[15:0];
    assign _1878 = { _1876, _1877 };
    assign _1886 = _1878 ^ _1885;
    assign _1887 = _1886[23:0];
    assign _1889 = { _1887, _1888 };
    assign _1904 = { _1889, _1903 };
    assign _1905 = _1904[511:64];
    assign _1922 = { _1905, _1920, _1921 };
    assign _1923 = _1922[511:224];
    assign _1934 = { _1923, _1932, _1933 };
    assign _1935 = _1934[511:384];
    assign _1937 = { _1935, _1928, _1936 };
    assign _1938 = _1937[511:416];
    assign _1940 = { _1938, _1927, _1939 };
    assign _1941 = _1940[511:96];
    assign _1958 = { _1941, _1956, _1957 };
    assign _1959 = _1958[511:256];
    assign _1970 = { _1959, _1968, _1969 };
    assign _1971 = _1970[511:288];
    assign _1973 = { _1971, _1964, _1972 };
    assign _1974 = _1973[511:448];
    assign _1976 = { _1974, _1963, _1975 };
    assign _1977 = _1976[511:128];
    assign _1994 = { _1977, _1992, _1993 };
    assign _1995 = _1994[511:160];
    assign _2006 = { _1995, _2004, _2005 };
    assign _2007 = _2006[511:320];
    assign _2009 = { _2007, _2000, _2008 };
    assign _2010 = _2009[511:480];
    assign _2012 = { _2010, _1999, _2011 };
    assign _2013 = _2012[511:32];
    assign _2029 = { _2013, _2028 };
    assign _2030 = _2029[511:160];
    assign _2041 = { _2030, _2039, _2040 };
    assign _2042 = _2041[511:288];
    assign _2044 = { _2042, _2035, _2043 };
    assign _2045 = _2044[511:416];
    assign _2047 = { _2045, _2034, _2046 };
    assign _2048 = _2047[511:64];
    assign _2065 = { _2048, _2063, _2064 };
    assign _2066 = _2065[511:192];
    assign _2077 = { _2066, _2075, _2076 };
    assign _2078 = _2077[511:320];
    assign _2080 = { _2078, _2071, _2079 };
    assign _2081 = _2080[511:448];
    assign _2083 = { _2081, _2070, _2082 };
    assign _2084 = _2083[511:96];
    assign _2101 = { _2084, _2099, _2100 };
    assign _2102 = _2101[511:224];
    assign _2113 = { _2102, _2111, _2112 };
    assign _2114 = _2113[511:352];
    assign _2116 = { _2114, _2107, _2115 };
    assign _2117 = _2116[511:480];
    assign _2119 = { _2117, _2106, _2118 };
    assign _2120 = _2119[511:480];
    assign _2124 = _2120 ^ _2123;
    assign _2125 = _2124[15:0];
    assign _2127 = { _2125, _2126 };
    assign _2135 = _2127 ^ _2134;
    assign _2136 = _2135[23:0];
    assign _2138 = { _2136, _2137 };
    assign _2154 = { _2138, _2153 };
    assign _2155 = _2154[511:480];
    assign _2159 = _2155 ^ _2158;
    assign _2160 = _2159[15:0];
    assign _2162 = { _2160, _2161 };
    assign _2170 = _2162 ^ _2169;
    assign _2171 = _2170[23:0];
    assign _2173 = { _2171, _2172 };
    assign _2188 = { _2173, _2187 };
    assign _2189 = _2188[511:64];
    assign _2206 = { _2189, _2204, _2205 };
    assign _2207 = _2206[511:224];
    assign _2218 = { _2207, _2216, _2217 };
    assign _2219 = _2218[511:384];
    assign _2221 = { _2219, _2212, _2220 };
    assign _2222 = _2221[511:416];
    assign _2224 = { _2222, _2211, _2223 };
    assign _2225 = _2224[511:96];
    assign _2242 = { _2225, _2240, _2241 };
    assign _2243 = _2242[511:256];
    assign _2254 = { _2243, _2252, _2253 };
    assign _2255 = _2254[511:288];
    assign _2257 = { _2255, _2248, _2256 };
    assign _2258 = _2257[511:448];
    assign _2260 = { _2258, _2247, _2259 };
    assign _2261 = _2260[511:128];
    assign _2278 = { _2261, _2276, _2277 };
    assign _2279 = _2278[511:160];
    assign _2290 = { _2279, _2288, _2289 };
    assign _2291 = _2290[511:320];
    assign _2293 = { _2291, _2284, _2292 };
    assign _2294 = _2293[511:480];
    assign _2296 = { _2294, _2283, _2295 };
    assign _2297 = _2296[511:32];
    assign _2313 = { _2297, _2312 };
    assign _2314 = _2313[511:160];
    assign _2325 = { _2314, _2323, _2324 };
    assign _2326 = _2325[511:288];
    assign _2328 = { _2326, _2319, _2327 };
    assign _2329 = _2328[511:416];
    assign _2331 = { _2329, _2318, _2330 };
    assign _2332 = _2331[511:64];
    assign _2349 = { _2332, _2347, _2348 };
    assign _2350 = _2349[511:192];
    assign _2361 = { _2350, _2359, _2360 };
    assign _2362 = _2361[511:320];
    assign _2364 = { _2362, _2355, _2363 };
    assign _2365 = _2364[511:448];
    assign _2367 = { _2365, _2354, _2366 };
    assign _2368 = _2367[511:96];
    assign _2385 = { _2368, _2383, _2384 };
    assign _2386 = _2385[511:224];
    assign _2397 = { _2386, _2395, _2396 };
    assign _2398 = _2397[511:352];
    assign _2400 = { _2398, _2391, _2399 };
    assign _2401 = _2400[511:480];
    assign _2403 = { _2401, _2390, _2402 };
    assign _2404 = _2403[511:480];
    assign _2408 = _2404 ^ _2407;
    assign _2409 = _2408[15:0];
    assign _2411 = { _2409, _2410 };
    assign _2419 = _2411 ^ _2418;
    assign _2420 = _2419[23:0];
    assign _2422 = { _2420, _2421 };
    assign _2438 = { _2422, _2437 };
    assign _2439 = _2438[511:480];
    assign _2443 = _2439 ^ _2442;
    assign _2444 = _2443[15:0];
    assign _2446 = { _2444, _2445 };
    assign _2454 = _2446 ^ _2453;
    assign _2455 = _2454[23:0];
    assign _2457 = { _2455, _2456 };
    assign _2472 = { _2457, _2471 };
    assign _2473 = _2472[511:64];
    assign _2490 = { _2473, _2488, _2489 };
    assign _2491 = _2490[511:224];
    assign _2502 = { _2491, _2500, _2501 };
    assign _2503 = _2502[511:384];
    assign _2505 = { _2503, _2496, _2504 };
    assign _2506 = _2505[511:416];
    assign _2508 = { _2506, _2495, _2507 };
    assign _2509 = _2508[511:96];
    assign _2526 = { _2509, _2524, _2525 };
    assign _2527 = _2526[511:256];
    assign _2538 = { _2527, _2536, _2537 };
    assign _2539 = _2538[511:288];
    assign _2541 = { _2539, _2532, _2540 };
    assign _2542 = _2541[511:448];
    assign _2544 = { _2542, _2531, _2543 };
    assign _2545 = _2544[511:128];
    assign _2562 = { _2545, _2560, _2561 };
    assign _2563 = _2562[511:160];
    assign _2574 = { _2563, _2572, _2573 };
    assign _2575 = _2574[511:320];
    assign _2577 = { _2575, _2568, _2576 };
    assign _2578 = _2577[511:480];
    assign _2580 = { _2578, _2567, _2579 };
    assign _2581 = _2580[511:32];
    assign _2597 = { _2581, _2596 };
    assign _2598 = _2597[511:160];
    assign _2609 = { _2598, _2607, _2608 };
    assign _2610 = _2609[511:288];
    assign _2612 = { _2610, _2603, _2611 };
    assign _2613 = _2612[511:416];
    assign _2615 = { _2613, _2602, _2614 };
    assign _2616 = _2615[511:64];
    assign _2633 = { _2616, _2631, _2632 };
    assign _2634 = _2633[511:192];
    assign _2645 = { _2634, _2643, _2644 };
    assign _2646 = _2645[511:320];
    assign _2648 = { _2646, _2639, _2647 };
    assign _2649 = _2648[511:448];
    assign _2651 = { _2649, _2638, _2650 };
    assign _2652 = _2651[511:96];
    assign _2669 = { _2652, _2667, _2668 };
    assign _2670 = _2669[511:224];
    assign _2681 = { _2670, _2679, _2680 };
    assign _2682 = _2681[511:352];
    assign _2684 = { _2682, _2675, _2683 };
    assign _2685 = _2684[511:480];
    assign _2687 = { _2685, _2674, _2686 };
    assign _2688 = _2687[511:480];
    assign _2692 = _2688 ^ _2691;
    assign _2693 = _2692[15:0];
    assign _2695 = { _2693, _2694 };
    assign _2703 = _2695 ^ _2702;
    assign _2704 = _2703[23:0];
    assign _2706 = { _2704, _2705 };
    assign _2722 = { _2706, _2721 };
    assign _2723 = _2722[511:480];
    assign _2727 = _2723 ^ _2726;
    assign _2728 = _2727[15:0];
    assign _2730 = { _2728, _2729 };
    assign _2738 = _2730 ^ _2737;
    assign _2739 = _2738[23:0];
    assign _2741 = { _2739, _2740 };
    assign _2756 = { _2741, _2755 };
    assign _2757 = _2756[511:64];
    assign _2774 = { _2757, _2772, _2773 };
    assign _2775 = _2774[511:224];
    assign _2786 = { _2775, _2784, _2785 };
    assign _2787 = _2786[511:384];
    assign _2789 = { _2787, _2780, _2788 };
    assign _2790 = _2789[511:416];
    assign _2792 = { _2790, _2779, _2791 };
    assign _2793 = _2792[511:96];
    assign _2810 = { _2793, _2808, _2809 };
    assign _2811 = _2810[511:256];
    assign _2822 = { _2811, _2820, _2821 };
    assign _2823 = _2822[511:288];
    assign _2825 = { _2823, _2816, _2824 };
    assign _2826 = _2825[511:448];
    assign _2828 = { _2826, _2815, _2827 };
    assign _2829 = _2828[511:128];
    assign _2846 = { _2829, _2844, _2845 };
    assign _2847 = _2846[511:160];
    assign _2858 = { _2847, _2856, _2857 };
    assign _2859 = _2858[511:320];
    assign _2861 = { _2859, _2852, _2860 };
    assign _2862 = _2861[511:480];
    assign _2864 = { _2862, _2851, _2863 };
    assign _2865 = _2864[511:480];
    assign _2 = clear;
    assign _4 = clock;
    assign _21 = _16[383:0];
    assign _18 = _16[415:384];
    assign _20 = _18 + _19;
    assign _17 = _16[511:416];
    assign _22 = { _17, _20, _21 };
    assign _6 = set_state;
    assign _12 = _6 == _11;
    assign _23 = _12 ? _9 : _22;
    assign _7 = _23;
    always @(posedge _4) begin
        if (_2)
            _16 <= _14;
        else
            _16 <= _7;
    end
    assign _24 = _16[511:480];
    assign _2866 = _24 + _2865;
    assign _2912 = { _2866, _2869, _2872, _2875, _2878, _2881, _2884, _2887, _2890, _2893, _2896, _2899, _2902, _2905, _2908, _2911 };
    assign _9 = round_input;
    assign _2913 = _9 ^ _2912;

    /* aliases */

    /* output assignments */
    assign round_output = _2913;

endmodule
