module poly1305_serial_encoder (
    clear,
    clock,
    number_of_input_bytes_minus_one,
    round_input,
    key,
    start,
    tag
);

    input clear;
    input clock;
    input [3:0] number_of_input_bytes_minus_one;
    input [127:0] round_input;
    input [255:0] key;
    input start;
    output [127:0] tag;

    /* signal declarations */
    wire [127:0] _95;
    wire vdd = 1'b1;
    wire [129:0] _46 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire _2;
    wire [129:0] _45 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire _4;
    wire [129:0] _92 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [258:0] _87 = 259'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011;
    wire [258:0] _81;
    wire [257:0] _82;
    wire _80 = 1'b0;
    wire [258:0] _83;
    wire [258:0] _75 = 259'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101;
    wire [517:0] _76;
    wire [258:0] _77;
    wire [258:0] _74 = 259'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [517:0] _78;
    wire [258:0] _79;
    wire [258:0] _84;
    wire [129:0] _85;
    wire [128:0] _73 = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [258:0] _86;
    wire [517:0] _88;
    wire [258:0] _89;
    wire [129:0] _67 = 130'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _66 = 130'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _65 = 130'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _64 = 130'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _63 = 130'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _62 = 130'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _61 = 130'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _60 = 130'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _59 = 130'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;
    wire [129:0] _58 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
    wire [129:0] _57 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
    wire [129:0] _56 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
    wire [129:0] _55 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;
    wire [129:0] _54 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
    wire [129:0] _53 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
    wire [129:0] _52 = 130'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
    wire [3:0] _6;
    reg [129:0] _68;
    wire [127:0] _8;
    wire [1:0] _50 = 2'b00;
    wire [129:0] _51;
    wire [129:0] _69;
    wire [130:0] _70;
    wire gnd = 1'b0;
    wire [130:0] _49;
    wire [130:0] _71;
    wire [7:0] _42;
    wire [7:0] _41;
    wire [7:0] _40;
    wire [7:0] _38;
    wire [7:0] _39;
    wire [7:0] _36;
    wire [7:0] _37;
    wire [7:0] _35;
    wire [7:0] _34;
    wire [7:0] _32;
    wire [7:0] _33;
    wire [7:0] _30;
    wire [7:0] _31;
    wire [7:0] _29;
    wire [7:0] _28;
    wire [7:0] _26;
    wire [7:0] _27;
    wire [7:0] _24 = 8'b11111100;
    wire [7:0] _23;
    wire [7:0] _25;
    wire [7:0] _22;
    wire [7:0] _21;
    wire [7:0] _19 = 8'b00001111;
    wire [255:0] _10;
    wire [127:0] _17;
    wire [7:0] _18;
    wire [7:0] _20;
    wire [127:0] _43;
    wire [258:0] _72;
    wire [258:0] _90;
    wire [129:0] _91;
    wire _15 = 1'b1;
    wire _12;
    wire _16;
    wire [129:0] _93;
    wire [129:0] _13;
    reg [129:0] _48;
    wire [127:0] _94;
    wire [127:0] _96;

    /* logic */
    assign _95 = _10[255:128];
    assign _2 = clear;
    assign _4 = clock;
    assign _81 = _72 - _79;
    assign _82 = _81[258:1];
    assign _83 = { _80, _82 };
    assign _76 = _72 * _75;
    assign _77 = _76[517:259];
    assign _78 = { _74, _77 };
    assign _79 = _78[258:0];
    assign _84 = _79 + _83;
    assign _85 = _84[258:129];
    assign _86 = { _73, _85 };
    assign _88 = _86 * _87;
    assign _89 = _88[258:0];
    assign _6 = number_of_input_bytes_minus_one;
    always @* begin
        case (_6)
        0: _68 <= _52;
        1: _68 <= _53;
        2: _68 <= _54;
        3: _68 <= _55;
        4: _68 <= _56;
        5: _68 <= _57;
        6: _68 <= _58;
        7: _68 <= _59;
        8: _68 <= _60;
        9: _68 <= _61;
        10: _68 <= _62;
        11: _68 <= _63;
        12: _68 <= _64;
        13: _68 <= _65;
        14: _68 <= _66;
        default: _68 <= _67;
        endcase
    end
    assign _8 = round_input;
    assign _51 = { _50, _8 };
    assign _69 = _51 | _68;
    assign _70 = { gnd, _69 };
    assign _49 = { gnd, _48 };
    assign _71 = _49 + _70;
    assign _42 = _17[7:0];
    assign _41 = _17[15:8];
    assign _40 = _17[23:16];
    assign _38 = _17[31:24];
    assign _39 = _38 & _19;
    assign _36 = _17[39:32];
    assign _37 = _36 & _24;
    assign _35 = _17[47:40];
    assign _34 = _17[55:48];
    assign _32 = _17[63:56];
    assign _33 = _32 & _19;
    assign _30 = _17[71:64];
    assign _31 = _30 & _24;
    assign _29 = _17[79:72];
    assign _28 = _17[87:80];
    assign _26 = _17[95:88];
    assign _27 = _26 & _19;
    assign _23 = _17[103:96];
    assign _25 = _23 & _24;
    assign _22 = _17[111:104];
    assign _21 = _17[119:112];
    assign _10 = key;
    assign _17 = _10[127:0];
    assign _18 = _17[127:120];
    assign _20 = _18 & _19;
    assign _43 = { _20, _21, _22, _25, _27, _28, _29, _31, _33, _34, _35, _37, _39, _40, _41, _42 };
    assign _72 = _43 * _71;
    assign _90 = _72 - _89;
    assign _91 = _90[129:0];
    assign _12 = start;
    assign _16 = _12 == _15;
    assign _93 = _16 ? _92 : _91;
    assign _13 = _93;
    always @(posedge _4) begin
        if (_2)
            _48 <= _46;
        else
            _48 <= _13;
    end
    assign _94 = _48[127:0];
    assign _96 = _94 + _95;

    /* aliases */

    /* output assignments */
    assign tag = _96;

endmodule
